
        library ieee;
        use ieee.std_logic_1164.all;
        use ieee.numeric_std.all;
        use ieee.std_logic_unsigned.all;

        entity project_tb is
        end project_tb;

        architecture projecttb of project_tb is
        constant c_CLOCK_PERIOD		: time := 100 ns;
        signal   tb_done		: std_logic;
        signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
        signal   tb_rst	                : std_logic := '0';
        signal   tb_start		: std_logic := '0';
        signal   tb_clk		        : std_logic := '0';
        signal   mem_o_data,mem_i_data	: std_logic_vector (7 downto 0);
        signal   enable_wire  		: std_logic;
        signal   mem_we		        : std_logic;

        type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
        type int_arr is array (0 to 1499) of integer range 0 to 255;
        shared variable addrs : int_arr :=(124, 111, 78, 46, 33, 83, 80, 59, 40, 51, 10, 54, 108, 106, 71, 40, 109, 89, 126, 3, 92, 44, 113, 120, 46, 9, 65, 90, 1, 15, 72, 8, 23, 123, 9, 16, 78, 7, 14, 49, 90, 15, 100, 5, 101, 78, 24, 115, 125, 65, 40, 60, 109, 106, 79, 18, 115, 81, 94, 84, 80, 73, 102, 35, 74, 33, 59, 16, 50, 8, 50, 100, 40, 97, 53, 127, 27, 11, 31, 102, 12, 72, 58, 82, 71, 101, 71, 117, 111, 114, 81, 64, 119, 62, 1, 65, 76, 28, 86, 123, 94, 20, 23, 10, 23, 97, 38, 75, 49, 116, 81, 9, 2, 44, 64, 103, 75, 88, 92, 50, 42, 93, 12, 69, 104, 27, 27, 38, 84, 77, 64, 50, 33, 112, 58, 95, 93, 125, 127, 32, 58, 90, 1, 23, 29, 2, 127, 28, 104, 29, 62, 20, 32, 48, 38, 85, 57, 31, 123, 123, 71, 120, 20, 59, 58, 53, 72, 88, 76, 121, 80, 12, 49, 105, 11, 3, 43, 64, 114, 23, 96, 47, 42, 28, 121, 4, 126, 14, 52, 85, 44, 4, 25, 24, 114, 24, 115, 80, 63, 78, 4, 65, 60, 89, 113, 49, 83, 49, 94, 19, 103, 14, 77, 64, 123, 3, 47, 97, 34, 23, 32, 8, 24, 37, 19, 21, 17, 116, 2, 43, 121, 51, 30, 31, 49, 121, 108, 110, 4, 92, 120, 118, 62, 105, 114, 107, 35, 64, 76, 37, 115, 121, 60, 55, 20, 56, 124, 87, 43, 36, 4, 107, 46, 45, 86, 33, 98, 17, 105, 12, 67, 86, 105, 50, 112, 82, 78, 69, 22, 10, 114, 111, 110, 95, 42, 71, 51, 81, 23, 32, 82, 49, 25, 47, 75, 35, 96, 100, 0, 28, 18, 72, 69, 109, 39, 18, 111, 69, 80, 91, 65, 78, 24, 46, 9, 117, 84, 75, 100, 105, 127, 20, 68, 111, 39, 50, 120, 38, 22, 15, 46, 45, 98, 107, 47, 84, 108, 28, 94, 55, 39, 79, 3, 105, 84, 96, 46, 65, 113, 78, 96, 113, 103, 108, 57, 1, 86, 34, 0, 10, 21, 69, 25, 40, 48, 92, 13, 77, 44, 109, 100, 44, 70, 36, 75, 116, 2, 61, 61, 58, 74, 33, 81, 63, 3, 14, 15, 122, 110, 67, 15, 19, 98, 60, 99, 54, 103, 30, 104, 48, 81, 44, 13, 33, 91, 126, 94, 53, 96, 69, 69, 81, 109, 59, 95, 13, 100, 116, 20, 54, 53, 101, 6, 6, 104, 47, 9, 51, 44, 6, 7, 9, 92, 76, 91, 114, 5, 92, 54, 32, 34, 72, 85, 3, 25, 51, 23, 92, 13, 46, 89, 87, 107, 78, 105, 19, 4, 63, 81, 28, 15, 109, 95, 85, 46, 69, 93, 74, 31, 119, 109, 16, 90, 43, 122, 18, 127, 87, 96, 65, 23, 11, 98, 30, 96, 35, 58, 112, 75, 73, 62, 56, 122, 106, 83, 103, 91, 19, 111, 79, 8, 94, 97, 47, 14, 38, 43, 56, 32, 47, 107, 10, 99, 97, 49, 112, 70, 122, 116, 107, 97, 112, 93, 0, 125, 89, 59, 19, 21, 59, 64, 39, 87, 115, 126, 40, 7, 8, 119, 98, 91, 106, 70, 109, 5, 51, 17, 121, 123, 100, 86, 46, 121, 34, 41, 31, 32, 3, 70, 124, 85, 46, 62, 85, 94, 69, 13, 127, 88, 13, 34, 92, 72, 4, 95, 126, 48, 43, 70, 10, 47, 39, 6, 23, 9, 30, 15, 66, 35, 51, 81, 95, 30, 42, 97, 2, 45, 80, 73, 36, 69, 61, 124, 14, 69, 43, 20, 52, 111, 101, 3, 120, 18, 40, 100, 38, 100, 0, 76, 120, 61, 61, 87, 48, 120, 85, 46, 15, 54, 97, 32, 3, 89, 16, 95, 5, 16, 82, 45, 55, 104, 8, 25, 108, 15, 40, 6, 53, 81, 23, 54, 112, 44, 48, 114, 9, 10, 113, 93, 2, 60, 24, 85, 125, 13, 49, 68, 4, 110, 89, 96, 63, 106, 99, 115, 28, 56, 30, 30, 47, 89, 1, 105, 92, 67, 60, 108, 71, 11, 11, 70, 53, 121, 1, 108, 117, 127, 82, 25, 8, 107, 36, 101, 105, 12, 110, 34, 10, 110, 51, 57, 97, 71, 99, 100, 85, 60, 90, 111, 114, 121, 55, 65, 27, 8, 40, 90, 4, 1, 72, 87, 12, 31, 26, 107, 3, 42, 2, 19, 88, 56, 89, 112, 22, 6, 102, 103, 51, 57, 54, 30, 2, 17, 109, 1, 32, 97, 78, 67, 46, 36, 22, 58, 72, 110, 124, 52, 119, 74, 16, 71, 28, 76, 24, 78, 112, 68, 3, 80, 65, 18, 62, 8, 35, 79, 41, 12, 76, 1, 59, 57, 72, 56, 120, 77, 16, 102, 29, 85, 50, 37, 29, 61, 92, 125, 116, 93, 122, 19, 99, 93, 90, 28, 66, 69, 47, 41, 23, 90, 103, 32, 28, 99, 23, 14, 8, 8, 60, 64, 38, 72, 127, 5, 23, 127, 48, 4, 40, 13, 102, 51, 71, 83, 23, 47, 40, 49, 28, 126, 57, 20, 122, 65, 16, 29, 53, 6, 6, 57, 123, 123, 28, 107, 25, 40, 4, 11, 39, 77, 76, 29, 52, 97, 96, 13, 95, 52, 79, 24, 52, 94, 119, 1, 87, 6, 29, 105, 18, 103, 100, 92, 79, 33, 59, 103, 117, 92, 115, 49, 107, 26, 92, 72, 54, 31, 37, 71, 16, 117, 36, 25, 97, 75, 94, 9, 110, 100, 109, 98, 83, 51, 25, 18, 106, 121, 81, 86, 66, 80, 124, 19, 120, 36, 41, 69, 112, 113, 56, 30, 46, 112, 72, 77, 25, 72, 58, 104, 24, 122, 97, 125, 3, 14, 100, 101, 41, 106, 24, 28, 68, 73, 91, 38, 1, 20, 21, 67, 2, 66, 51, 10, 56, 119, 89, 46, 16, 18, 103, 46, 24, 116, 26, 12, 50, 43, 81, 9, 61, 94, 104, 18, 29, 103, 22, 91, 88, 13, 44, 35, 0, 76, 82, 16, 66, 75, 127, 65, 126, 118, 99, 9, 39, 19, 54, 59, 50, 35, 65, 46, 33, 74, 86, 107, 37, 49, 122, 32, 47, 76, 103, 41, 62, 12, 48, 109, 98, 25, 51, 72, 110, 79, 90, 73, 118, 63, 66, 5, 22, 120, 98, 80, 16, 18, 7, 49, 13, 96, 54, 44, 25, 68, 86, 1, 91, 74, 18, 12, 100, 40, 102, 92, 62, 9, 65, 121, 35, 25, 3, 40, 32, 85, 110, 88, 3, 115, 107, 107, 114, 48, 2, 92, 57, 121, 122, 41, 53, 96, 22, 113, 10, 65, 42, 119, 123, 119, 71, 100, 2, 108, 84, 1, 119, 13, 126, 90, 26, 25, 52, 11, 12, 90, 44, 53, 58, 65, 3, 83, 10, 91, 65, 9, 95, 15, 12, 33, 74, 0, 125, 78, 88, 67, 78, 18, 64, 35, 57, 114, 9, 83, 16, 124, 34, 58, 27, 95, 109, 8, 60, 31, 54, 98, 67, 113, 112, 36, 29, 100, 77, 82, 127, 10, 60, 19, 18, 3, 30, 124, 46, 104, 29, 95, 65, 83, 8, 19, 58, 124, 84, 14, 119, 69, 50, 1, 2, 10, 93, 120, 17, 18, 101, 112, 15, 26, 82, 59, 110, 98, 78, 91, 108, 72, 15, 71, 8, 21, 43, 79, 51, 31, 38, 54, 31, 83, 76, 55, 73, 104, 84, 16, 93, 61, 16, 112, 27, 68, 38, 55, 34, 85, 53, 51, 123, 5, 78, 120, 60, 102, 109, 69, 102, 86, 81, 38, 16, 100, 104, 85, 38, 60, 119, 43, 64, 109, 121, 2, 57, 68, 21, 116, 121, 90, 68, 10, 23, 4, 3, 110, 23, 26, 71, 113, 98, 85, 93, 84, 73, 113, 95, 117, 42, 39, 2, 66, 83, 27, 41, 33, 51, 6, 19, 107, 10, 32, 81, 112, 16, 91, 38, 0, 80, 96, 55, 44, 49, 59, 59, 127, 14, 22, 104, 111, 41, 106, 82, 111, 18, 79, 65, 104, 34, 1, 83, 16, 20, 79, 93, 112, 97, 58, 90, 28, 107, 104, 89, 127, 27, 8, 107, 10, 127, 56, 43, 49, 99, 105, 85, 84, 38, 69, 34, 5, 10, 98, 13, 83, 64, 120, 27, 103, 40, 114, 11, 109, 124, 94, 51, 41, 96, 111, 26, 47, 71, 70, 103, 65, 37, 71, 90, 77, 31, 54, 110, 124, 36, 70, 13, 116, 61, 22, 117, 36, 51, 11, 19, 70, 113, 13, 100, 81, 15, 95, 24, 18, 113, 77, 122, 3, 28, 104, 104, 42, 103, 119, 39, 126, 63, 5, 71, 80, 25, 79, 101, 110, 111, 11, 104, 90, 92, 21, 77, 99, 13, 27, 33, 19, 117, 24, 20, 111, 9, 24, 60, 63, 53, 63, 47, 102, 71, 59, 103, 91, 3, 16, 75, 47, 68, 71, 112, 23, 12, 102, 29, 116, 92, 55, 67, 1, 34, 69, 57, 20, 111, 61, 90, 41, 38, 49, 41, 114, 109, 74, 0, 92, 69, 24, 70, 97, 59, 23, 40);
shared variable enc_addrs : int_arr :=(232, 111, 78, 248, 145, 83, 80, 209, 148, 51, 10, 54, 108, 106, 71, 40, 109, 89, 126, 3, 241, 44, 113, 145, 46, 9, 65, 90, 1, 161, 72, 8, 23, 123, 132, 16, 78, 7, 168, 49, 90, 15, 100, 5, 101, 78, 24, 115, 125, 193, 40, 60, 109, 106, 79, 18, 115, 81, 178, 84, 80, 73, 102, 209, 74, 33, 178, 16, 50, 129, 216, 100, 40, 168, 53, 127, 27, 11, 31, 193, 12, 72, 58, 82, 162, 101, 71, 117, 111, 114, 81, 161, 119, 62, 1, 65, 225, 196, 232, 123, 232, 20, 228, 10, 178, 145, 38, 75, 49, 116, 145, 9, 2, 44, 193, 103, 161, 88, 92, 50, 42, 93, 12, 69, 104, 210, 228, 248, 129, 177, 64, 50, 33, 112, 58, 95, 93, 125, 127, 32, 58, 90, 209, 193, 29, 2, 127, 196, 104, 168, 62, 194, 32, 48, 38, 85, 164, 31, 123, 194, 71, 120, 20, 164, 58, 53, 216, 212, 76, 121, 80, 12, 49, 105, 130, 3, 43, 196, 114, 145, 96, 47, 42, 28, 121, 4, 126, 14, 52, 232, 44, 209, 25, 24, 114, 24, 115, 209, 63, 244, 4, 65, 60, 145, 113, 49, 83, 49, 94, 145, 103, 168, 77, 64, 161, 3, 148, 97, 34, 23, 32, 8, 168, 37, 19, 21, 145, 116, 2, 43, 121, 51, 30, 161, 49, 121, 108, 194, 4, 92, 120, 118, 62, 161, 114, 184, 35, 64, 76, 37, 115, 121, 60, 55, 20, 56, 124, 225, 43, 36, 4, 193, 46, 210, 86, 130, 98, 17, 105, 129, 67, 86, 105, 50, 216, 82, 78, 152, 210, 10, 114, 111, 110, 95, 42, 71, 51, 81, 23, 161, 82, 168, 25, 47, 75, 35, 96, 132, 0, 28, 209, 226, 69, 130, 39, 226, 111, 69, 80, 91, 212, 78, 196, 46, 9, 117, 84, 168, 100, 105, 127, 20, 68, 111, 226, 162, 120, 145, 22, 226, 46, 45, 98, 107, 216, 84, 178, 28, 94, 55, 226, 79, 3, 162, 84, 136, 46, 65, 113, 78, 196, 194, 103, 108, 57, 1, 86, 241, 0, 146, 21, 69, 200, 232, 48, 92, 13, 77, 44, 168, 216, 44, 212, 248, 178, 145, 196, 61, 196, 216, 74, 33, 81, 63, 193, 14, 15, 122, 110, 67, 193, 19, 130, 60, 99, 184, 103, 30, 104, 164, 81, 148, 13, 162, 91, 126, 94, 53, 96, 69, 69, 81, 109, 59, 95, 13, 225, 116, 20, 184, 53, 101, 6, 6, 104, 47, 9, 51, 44, 241, 242, 9, 180, 76, 91, 114, 5, 92, 54, 216, 34, 72, 164, 3, 25, 51, 23, 196, 13, 46, 145, 200, 107, 164, 242, 19, 4, 130, 180, 28, 15, 109, 225, 85, 46, 69, 93, 74, 226, 119, 109, 16, 90, 152, 122, 18, 127, 168, 96, 225, 210, 11, 98, 196, 96, 35, 58, 112, 75, 152, 62, 130, 122, 106, 83, 103, 216, 241, 111, 79, 8, 94, 97, 47, 14, 38, 228, 130, 209, 47, 193, 130, 99, 97, 49, 216, 70, 122, 145, 107, 97, 212, 93, 0, 125, 193, 59, 130, 21, 152, 64, 39, 87, 115, 126, 40, 7, 8, 119, 98, 91, 184, 70, 109, 5, 51, 17, 121, 123, 184, 148, 148, 244, 34, 41, 31, 32, 180, 70, 124, 85, 46, 62, 85, 94, 69, 13, 127, 88, 13, 34, 92, 72, 4, 95, 126, 48, 43, 216, 10, 47, 39, 6, 23, 148, 30, 177, 209, 35, 51, 180, 95, 30, 42, 161, 2, 178, 80, 228, 36, 69, 129, 124, 14, 69, 43, 20, 52, 111, 101, 3, 120, 18, 40, 100, 194, 100, 129, 76, 210, 61, 61, 226, 48, 194, 85, 46, 15, 178, 97, 32, 3, 89, 16, 95, 5, 16, 180, 177, 55, 104, 244, 25, 108, 15, 136, 178, 248, 212, 129, 54, 112, 44, 164, 114, 9, 10, 146, 196, 177, 244, 193, 85, 125, 13, 49, 68, 4, 244, 89, 96, 196, 106, 99, 115, 28, 216, 30, 30, 152, 89, 1, 105, 92, 67, 242, 108, 71, 11, 11, 70, 53, 196, 1, 108, 117, 127, 132, 25, 8, 107, 36, 101, 105, 225, 110, 34, 10, 110, 232, 148, 97, 146, 99, 152, 85, 60, 90, 244, 114, 121, 55, 212, 27, 8, 209, 136, 4, 194, 72, 248, 244, 31, 26, 107, 3, 42, 226, 19, 88, 56, 89, 177, 22, 212, 102, 103, 136, 57, 146, 30, 2, 17, 109, 1, 32, 228, 78, 209, 46, 177, 161, 58, 72, 110, 130, 52, 146, 146, 16, 193, 28, 132, 148, 78, 112, 68, 145, 80, 132, 18, 62, 8, 35, 162, 41, 12, 161, 1, 59, 57, 72, 56, 120, 77, 16, 102, 29, 85, 50, 37, 29, 200, 92, 125, 116, 93, 122, 19, 99, 93, 90, 136, 66, 69, 136, 241, 184, 90, 180, 32, 28, 241, 23, 14, 8, 8, 228, 228, 38, 161, 127, 5, 23, 127, 146, 148, 40, 13, 102, 148, 71, 83, 23, 47, 226, 49, 28, 126, 57, 20, 122, 65, 209, 193, 53, 6, 6, 57, 123, 123, 194, 107, 25, 216, 4, 11, 39, 77, 148, 29, 52, 97, 96, 13, 95, 148, 79, 177, 52, 94, 119, 1, 87, 6, 178, 105, 18, 103, 100, 92, 79, 33, 59, 103, 117, 92, 177, 161, 241, 26, 92, 72, 54, 209, 37, 71, 16, 117, 36, 196, 184, 75, 242, 9, 110, 164, 109, 194, 83, 130, 25, 18, 106, 121, 81, 152, 66, 80, 124, 19, 193, 36, 41, 184, 112, 113, 56, 209, 193, 112, 72, 77, 25, 72, 58, 241, 209, 122, 97, 125, 3, 14, 100, 101, 41, 106, 24, 28, 68, 164, 146, 38, 145, 20, 145, 177, 2, 66, 51, 10, 56, 119, 89, 46, 180, 18, 226, 46, 24, 116, 161, 12, 50, 43, 216, 9, 129, 94, 216, 18, 29, 103, 22, 91, 88, 13, 44, 216, 0, 216, 228, 162, 242, 75, 127, 65, 126, 118, 99, 9, 39, 194, 54, 59, 50, 35, 65, 46, 33, 74, 86, 107, 37, 49, 122, 32, 47, 76, 193, 148, 162, 12, 48, 146, 98, 25, 51, 72, 110, 79, 90, 73, 118, 63, 66, 5, 244, 120, 98, 164, 16, 18, 148, 49, 13, 96, 178, 44, 25, 68, 86, 1, 91, 74, 18, 12, 100, 212, 102, 92, 216, 9, 65, 121, 35, 25, 3, 40, 32, 145, 110, 88, 3, 242, 242, 107, 114, 48, 2, 92, 57, 121, 122, 146, 53, 96, 130, 113, 162, 232, 226, 119, 123, 119, 71, 225, 161, 228, 248, 1, 216, 196, 126, 178, 26, 25, 52, 11, 12, 90, 44, 53, 58, 65, 3, 83, 200, 91, 65, 152, 225, 15, 12, 33, 74, 0, 125, 129, 88, 67, 78, 18, 64, 35, 57, 228, 132, 83, 16, 124, 34, 212, 27, 95, 109, 8, 60, 31, 193, 168, 209, 113, 112, 129, 29, 100, 77, 82, 127, 10, 196, 19, 18, 3, 30, 124, 46, 104, 132, 95, 65, 83, 248, 19, 132, 241, 84, 14, 119, 69, 248, 1, 2, 168, 152, 146, 17, 18, 101, 161, 15, 212, 148, 59, 110, 136, 162, 228, 108, 178, 132, 71, 8, 21, 43, 164, 51, 146, 38, 200, 31, 83, 76, 55, 73, 232, 84, 16, 161, 61, 16, 112, 27, 168, 180, 55, 34, 85, 53, 51, 123, 5, 78, 226, 60, 102, 242, 69, 102, 86, 81, 38, 16, 100, 104, 164, 38, 60, 119, 43, 64, 109, 121, 2, 57, 164, 21, 116, 121, 209, 68, 10, 196, 212, 3, 110, 23, 26, 71, 113, 98, 85, 148, 210, 73, 113, 95, 194, 42, 184, 2, 66, 83, 27, 41, 130, 51, 178, 161, 107, 10, 32, 81, 112, 16, 91, 38, 0, 228, 96, 55, 44, 130, 59, 59, 127, 14, 22, 180, 111, 41, 241, 82, 111, 18, 79, 65, 232, 34, 1, 83, 177, 20, 79, 93, 112, 97, 58, 148, 130, 107, 104, 209, 127, 27, 8, 107, 136, 127, 244, 43, 248, 99, 105, 145, 84, 38, 164, 164, 194, 10, 98, 13, 83, 64, 180, 27, 103, 40, 114, 11, 225, 124, 94, 51, 41, 129, 111, 26, 177, 71, 244, 194, 65, 37, 71, 90, 77, 136, 54, 110, 124, 36, 70, 13, 116, 161, 212, 117, 168, 51, 194, 19, 200, 113, 232, 100, 129, 15, 184, 148, 18, 113, 77, 130, 3, 28, 104, 241, 42, 103, 119, 39, 126, 63, 5, 71, 80, 25, 79, 216, 161, 111, 11, 104, 90, 209, 21, 77, 99, 178, 27, 33, 19, 117, 24, 20, 111, 248, 24, 60, 210, 53, 242, 47, 102, 136, 59, 129, 91, 232, 242, 200, 47, 68, 71, 112, 23, 12, 102, 194, 116, 92, 55, 67, 1, 34, 69, 57, 20, 111, 164, 90, 41, 38, 49, 130, 114, 200, 74, 0, 92, 168, 232, 70, 97, 59, 23, 40);

shared variable i : integer range 0 to 1501 := 0;
shared variable is_next : integer range 0 to 3 := 0;

-- come da esempio su specifica
signal RAM: ram_type := (0 => std_logic_vector(to_unsigned(43 , 8)),
                        1 => std_logic_vector(to_unsigned( 69 , 8)),
                        2 => std_logic_vector(to_unsigned( 0 , 8)),
                        3 => std_logic_vector(to_unsigned( 22 , 8)),
                        4 => std_logic_vector(to_unsigned( 35 , 8)),
                        5 => std_logic_vector(to_unsigned( 98 , 8)),
                        6 => std_logic_vector(to_unsigned( 121 , 8)),
                        7 => std_logic_vector(to_unsigned( 89 , 8)),
                        8 => std_logic_vector(to_unsigned( 124 , 8)),
            others => (others =>'0'));

component project_reti_logiche is
port (
    i_clk         : in  std_logic;
    i_start       : in  std_logic;
    i_rst         : in  std_logic;
    i_data        : in  std_logic_vector(7 downto 0);
    o_address     : out std_logic_vector(15 downto 0);
    o_done        : out std_logic;
    o_en          : out std_logic;
    o_we          : out std_logic;
    o_data        : out std_logic_vector (7 downto 0)
    );
end component project_reti_logiche;


begin
UUT: project_reti_logiche
port map (
        i_clk      	=> tb_clk,
        i_start       => tb_start,
        i_rst      	=> tb_rst,
        i_data    	=> mem_o_data,
        o_address  	=> mem_address,
        o_done      	=> tb_done,
        o_en   	=> enable_wire,
        o_we 		=> mem_we,
        o_data    	=> mem_i_data
        );

p_CLK_GEN : process is
begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
end process p_CLK_GEN;


MEM : process(tb_clk)
begin
    if tb_clk'event and tb_clk = '1' then
        if enable_wire = '1' then
            if mem_we = '1' then
                RAM(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 1 ns;
            else
                mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
            end if;
        end if;

         if i=1 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 121 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=2 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 59 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 108 , 8)),
                    4 => std_logic_vector(to_unsigned( 5 , 8)),
                    5 => std_logic_vector(to_unsigned( 91 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 104 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=3 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 33 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 21 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 124 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=4 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 33 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 21 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 124 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=5 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 31 , 8)),
                    2 => std_logic_vector(to_unsigned( 60 , 8)),
                    3 => std_logic_vector(to_unsigned( 104 , 8)),
                    4 => std_logic_vector(to_unsigned( 12 , 8)),
                    5 => std_logic_vector(to_unsigned( 8 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=6 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 16 , 8)),
                    2 => std_logic_vector(to_unsigned( 22 , 8)),
                    3 => std_logic_vector(to_unsigned( 26 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 12 , 8)),
                    7 => std_logic_vector(to_unsigned( 37 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=7 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 16 , 8)),
                    2 => std_logic_vector(to_unsigned( 22 , 8)),
                    3 => std_logic_vector(to_unsigned( 26 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 12 , 8)),
                    7 => std_logic_vector(to_unsigned( 37 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=8 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),
                    1 => std_logic_vector(to_unsigned( 38 , 8)),
                    2 => std_logic_vector(to_unsigned( 29 , 8)),
                    3 => std_logic_vector(to_unsigned( 57 , 8)),
                    4 => std_logic_vector(to_unsigned( 68 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 12 , 8)),
                    7 => std_logic_vector(to_unsigned( 64 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=9 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),
                    1 => std_logic_vector(to_unsigned( 108 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 65 , 8)),
                    4 => std_logic_vector(to_unsigned( 115 , 8)),
                    5 => std_logic_vector(to_unsigned( 99 , 8)),
                    6 => std_logic_vector(to_unsigned( 93 , 8)),
                    7 => std_logic_vector(to_unsigned( 55 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=10 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),
                    1 => std_logic_vector(to_unsigned( 108 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 65 , 8)),
                    4 => std_logic_vector(to_unsigned( 115 , 8)),
                    5 => std_logic_vector(to_unsigned( 99 , 8)),
                    6 => std_logic_vector(to_unsigned( 93 , 8)),
                    7 => std_logic_vector(to_unsigned( 55 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=11 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),
                    1 => std_logic_vector(to_unsigned( 17 , 8)),
                    2 => std_logic_vector(to_unsigned( 94 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 8 , 8)),
                    5 => std_logic_vector(to_unsigned( 3 , 8)),
                    6 => std_logic_vector(to_unsigned( 27 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=12 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 50 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 119 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 21 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=13 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 50 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 119 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 21 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=14 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 81 , 8)),
                    3 => std_logic_vector(to_unsigned( 3 , 8)),
                    4 => std_logic_vector(to_unsigned( 30 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 66 , 8)),
                    7 => std_logic_vector(to_unsigned( 55 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=15 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),
                    1 => std_logic_vector(to_unsigned( 14 , 8)),
                    2 => std_logic_vector(to_unsigned( 89 , 8)),
                    3 => std_logic_vector(to_unsigned( 28 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 122 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 9 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=16 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),
                    1 => std_logic_vector(to_unsigned( 14 , 8)),
                    2 => std_logic_vector(to_unsigned( 89 , 8)),
                    3 => std_logic_vector(to_unsigned( 28 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 122 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 9 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=17 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 26 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 54 , 8)),
                    6 => std_logic_vector(to_unsigned( 64 , 8)),
                    7 => std_logic_vector(to_unsigned( 96 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=18 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 34 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 66 , 8)),
                    5 => std_logic_vector(to_unsigned( 48 , 8)),
                    6 => std_logic_vector(to_unsigned( 60 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=19 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 34 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 66 , 8)),
                    5 => std_logic_vector(to_unsigned( 48 , 8)),
                    6 => std_logic_vector(to_unsigned( 60 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=20 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 99 , 8)),
                    2 => std_logic_vector(to_unsigned( 29 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 67 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 115 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=21 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 83, 8)),
                    1 => std_logic_vector(to_unsigned( 108 , 8)),
                    2 => std_logic_vector(to_unsigned( 23 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 66 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=22 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 83, 8)),
                    1 => std_logic_vector(to_unsigned( 108 , 8)),
                    2 => std_logic_vector(to_unsigned( 23 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 66 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=23 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 120 , 8)),
                    2 => std_logic_vector(to_unsigned( 104 , 8)),
                    3 => std_logic_vector(to_unsigned( 21 , 8)),
                    4 => std_logic_vector(to_unsigned( 73 , 8)),
                    5 => std_logic_vector(to_unsigned( 1 , 8)),
                    6 => std_logic_vector(to_unsigned( 111 , 8)),
                    7 => std_logic_vector(to_unsigned( 100 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=24 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 111 , 8)),
                    2 => std_logic_vector(to_unsigned( 78 , 8)),
                    3 => std_logic_vector(to_unsigned( 40 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 50 , 8)),
                    6 => std_logic_vector(to_unsigned( 28 , 8)),
                    7 => std_logic_vector(to_unsigned( 17 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=25 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 111 , 8)),
                    2 => std_logic_vector(to_unsigned( 78 , 8)),
                    3 => std_logic_vector(to_unsigned( 40 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 50 , 8)),
                    6 => std_logic_vector(to_unsigned( 28 , 8)),
                    7 => std_logic_vector(to_unsigned( 17 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=26 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 37 , 8)),
                    4 => std_logic_vector(to_unsigned( 8 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 120 , 8)),
                    7 => std_logic_vector(to_unsigned( 58 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=27 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 80, 8)),
                    1 => std_logic_vector(to_unsigned( 14 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 27 , 8)),
                    5 => std_logic_vector(to_unsigned( 7 , 8)),
                    6 => std_logic_vector(to_unsigned( 18 , 8)),
                    7 => std_logic_vector(to_unsigned( 59 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=28 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 80, 8)),
                    1 => std_logic_vector(to_unsigned( 14 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 27 , 8)),
                    5 => std_logic_vector(to_unsigned( 7 , 8)),
                    6 => std_logic_vector(to_unsigned( 18 , 8)),
                    7 => std_logic_vector(to_unsigned( 59 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=29 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 76, 8)),
                    1 => std_logic_vector(to_unsigned( 32 , 8)),
                    2 => std_logic_vector(to_unsigned( 15 , 8)),
                    3 => std_logic_vector(to_unsigned( 111 , 8)),
                    4 => std_logic_vector(to_unsigned( 20 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 105 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=30 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 4, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 13 , 8)),
                    3 => std_logic_vector(to_unsigned( 83 , 8)),
                    4 => std_logic_vector(to_unsigned( 55 , 8)),
                    5 => std_logic_vector(to_unsigned( 78 , 8)),
                    6 => std_logic_vector(to_unsigned( 48 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=31 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 4, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 13 , 8)),
                    3 => std_logic_vector(to_unsigned( 83 , 8)),
                    4 => std_logic_vector(to_unsigned( 55 , 8)),
                    5 => std_logic_vector(to_unsigned( 78 , 8)),
                    6 => std_logic_vector(to_unsigned( 48 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=32 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 88, 8)),
                    1 => std_logic_vector(to_unsigned( 120 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 7 , 8)),
                    5 => std_logic_vector(to_unsigned( 17 , 8)),
                    6 => std_logic_vector(to_unsigned( 65 , 8)),
                    7 => std_logic_vector(to_unsigned( 45 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=33 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),
                    1 => std_logic_vector(to_unsigned( 27 , 8)),
                    2 => std_logic_vector(to_unsigned( 50 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 13 , 8)),
                    5 => std_logic_vector(to_unsigned( 75 , 8)),
                    6 => std_logic_vector(to_unsigned( 31 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=34 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),
                    1 => std_logic_vector(to_unsigned( 27 , 8)),
                    2 => std_logic_vector(to_unsigned( 50 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 13 , 8)),
                    5 => std_logic_vector(to_unsigned( 75 , 8)),
                    6 => std_logic_vector(to_unsigned( 31 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=35 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 120 , 8)),
                    2 => std_logic_vector(to_unsigned( 100 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 82 , 8)),
                    5 => std_logic_vector(to_unsigned( 28 , 8)),
                    6 => std_logic_vector(to_unsigned( 70 , 8)),
                    7 => std_logic_vector(to_unsigned( 4 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=36 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 92 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 73 , 8)),
                    6 => std_logic_vector(to_unsigned( 14 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=37 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 92 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 73 , 8)),
                    6 => std_logic_vector(to_unsigned( 14 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=38 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 83, 8)),
                    1 => std_logic_vector(to_unsigned( 57 , 8)),
                    2 => std_logic_vector(to_unsigned( 11 , 8)),
                    3 => std_logic_vector(to_unsigned( 119 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 34 , 8)),
                    6 => std_logic_vector(to_unsigned( 109 , 8)),
                    7 => std_logic_vector(to_unsigned( 22 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=39 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 57 , 8)),
                    2 => std_logic_vector(to_unsigned( 53 , 8)),
                    3 => std_logic_vector(to_unsigned( 110 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 7 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 38 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=40 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 57 , 8)),
                    2 => std_logic_vector(to_unsigned( 53 , 8)),
                    3 => std_logic_vector(to_unsigned( 110 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 7 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 38 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=41 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 81, 8)),
                    1 => std_logic_vector(to_unsigned( 50 , 8)),
                    2 => std_logic_vector(to_unsigned( 117 , 8)),
                    3 => std_logic_vector(to_unsigned( 99 , 8)),
                    4 => std_logic_vector(to_unsigned( 10 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 23 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=42 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 33, 8)),
                    1 => std_logic_vector(to_unsigned( 107 , 8)),
                    2 => std_logic_vector(to_unsigned( 83 , 8)),
                    3 => std_logic_vector(to_unsigned( 39 , 8)),
                    4 => std_logic_vector(to_unsigned( 91 , 8)),
                    5 => std_logic_vector(to_unsigned( 8 , 8)),
                    6 => std_logic_vector(to_unsigned( 58 , 8)),
                    7 => std_logic_vector(to_unsigned( 1 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=43 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 33, 8)),
                    1 => std_logic_vector(to_unsigned( 107 , 8)),
                    2 => std_logic_vector(to_unsigned( 83 , 8)),
                    3 => std_logic_vector(to_unsigned( 39 , 8)),
                    4 => std_logic_vector(to_unsigned( 91 , 8)),
                    5 => std_logic_vector(to_unsigned( 8 , 8)),
                    6 => std_logic_vector(to_unsigned( 58 , 8)),
                    7 => std_logic_vector(to_unsigned( 1 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=44 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),
                    1 => std_logic_vector(to_unsigned( 84 , 8)),
                    2 => std_logic_vector(to_unsigned( 6 , 8)),
                    3 => std_logic_vector(to_unsigned( 66 , 8)),
                    4 => std_logic_vector(to_unsigned( 70 , 8)),
                    5 => std_logic_vector(to_unsigned( 115 , 8)),
                    6 => std_logic_vector(to_unsigned( 79 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=45 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),
                    1 => std_logic_vector(to_unsigned( 120 , 8)),
                    2 => std_logic_vector(to_unsigned( 65 , 8)),
                    3 => std_logic_vector(to_unsigned( 11 , 8)),
                    4 => std_logic_vector(to_unsigned( 39 , 8)),
                    5 => std_logic_vector(to_unsigned( 5 , 8)),
                    6 => std_logic_vector(to_unsigned( 52 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=46 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),
                    1 => std_logic_vector(to_unsigned( 120 , 8)),
                    2 => std_logic_vector(to_unsigned( 65 , 8)),
                    3 => std_logic_vector(to_unsigned( 11 , 8)),
                    4 => std_logic_vector(to_unsigned( 39 , 8)),
                    5 => std_logic_vector(to_unsigned( 5 , 8)),
                    6 => std_logic_vector(to_unsigned( 52 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=47 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),
                    1 => std_logic_vector(to_unsigned( 77 , 8)),
                    2 => std_logic_vector(to_unsigned( 98 , 8)),
                    3 => std_logic_vector(to_unsigned( 44 , 8)),
                    4 => std_logic_vector(to_unsigned( 60 , 8)),
                    5 => std_logic_vector(to_unsigned( 94 , 8)),
                    6 => std_logic_vector(to_unsigned( 120 , 8)),
                    7 => std_logic_vector(to_unsigned( 9 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=48 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 39, 8)),
                    1 => std_logic_vector(to_unsigned( 19 , 8)),
                    2 => std_logic_vector(to_unsigned( 27 , 8)),
                    3 => std_logic_vector(to_unsigned( 5 , 8)),
                    4 => std_logic_vector(to_unsigned( 65 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 77 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=49 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 39, 8)),
                    1 => std_logic_vector(to_unsigned( 19 , 8)),
                    2 => std_logic_vector(to_unsigned( 27 , 8)),
                    3 => std_logic_vector(to_unsigned( 5 , 8)),
                    4 => std_logic_vector(to_unsigned( 65 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 77 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=50 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 93 , 8)),
                    3 => std_logic_vector(to_unsigned( 31 , 8)),
                    4 => std_logic_vector(to_unsigned( 22 , 8)),
                    5 => std_logic_vector(to_unsigned( 77 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 118 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=51 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),
                    1 => std_logic_vector(to_unsigned( 114 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 87 , 8)),
                    5 => std_logic_vector(to_unsigned( 74 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 17 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=52 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),
                    1 => std_logic_vector(to_unsigned( 114 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 87 , 8)),
                    5 => std_logic_vector(to_unsigned( 74 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 17 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=53 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 68 , 8)),
                    3 => std_logic_vector(to_unsigned( 99 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 5 , 8)),
                    7 => std_logic_vector(to_unsigned( 12 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=54 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 42 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 34 , 8)),
                    6 => std_logic_vector(to_unsigned( 121 , 8)),
                    7 => std_logic_vector(to_unsigned( 20 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=55 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 42 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 34 , 8)),
                    6 => std_logic_vector(to_unsigned( 121 , 8)),
                    7 => std_logic_vector(to_unsigned( 20 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=56 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 62 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 67 , 8)),
                    5 => std_logic_vector(to_unsigned( 25 , 8)),
                    6 => std_logic_vector(to_unsigned( 31 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=57 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 20 , 8)),
                    3 => std_logic_vector(to_unsigned( 93 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 69 , 8)),
                    7 => std_logic_vector(to_unsigned( 107 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=58 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 20 , 8)),
                    3 => std_logic_vector(to_unsigned( 93 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 69 , 8)),
                    7 => std_logic_vector(to_unsigned( 107 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=59 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 77, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 114 , 8)),
                    3 => std_logic_vector(to_unsigned( 40 , 8)),
                    4 => std_logic_vector(to_unsigned( 3 , 8)),
                    5 => std_logic_vector(to_unsigned( 73 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 108 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=60 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 12 , 8)),
                    3 => std_logic_vector(to_unsigned( 66 , 8)),
                    4 => std_logic_vector(to_unsigned( 22 , 8)),
                    5 => std_logic_vector(to_unsigned( 37 , 8)),
                    6 => std_logic_vector(to_unsigned( 7 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=61 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 12 , 8)),
                    3 => std_logic_vector(to_unsigned( 66 , 8)),
                    4 => std_logic_vector(to_unsigned( 22 , 8)),
                    5 => std_logic_vector(to_unsigned( 37 , 8)),
                    6 => std_logic_vector(to_unsigned( 7 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=62 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 47, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 64 , 8)),
                    3 => std_logic_vector(to_unsigned( 3 , 8)),
                    4 => std_logic_vector(to_unsigned( 33 , 8)),
                    5 => std_logic_vector(to_unsigned( 25 , 8)),
                    6 => std_logic_vector(to_unsigned( 59 , 8)),
                    7 => std_logic_vector(to_unsigned( 39 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=63 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),
                    1 => std_logic_vector(to_unsigned( 2 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 45 , 8)),
                    4 => std_logic_vector(to_unsigned( 124 , 8)),
                    5 => std_logic_vector(to_unsigned( 35 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 19 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=64 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),
                    1 => std_logic_vector(to_unsigned( 2 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 45 , 8)),
                    4 => std_logic_vector(to_unsigned( 124 , 8)),
                    5 => std_logic_vector(to_unsigned( 35 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 19 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=65 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 27 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 98 , 8)),
                    4 => std_logic_vector(to_unsigned( 92 , 8)),
                    5 => std_logic_vector(to_unsigned( 0 , 8)),
                    6 => std_logic_vector(to_unsigned( 88 , 8)),
                    7 => std_logic_vector(to_unsigned( 37 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=66 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 48 , 8)),
                    2 => std_logic_vector(to_unsigned( 12 , 8)),
                    3 => std_logic_vector(to_unsigned( 58 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=67 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 48 , 8)),
                    2 => std_logic_vector(to_unsigned( 12 , 8)),
                    3 => std_logic_vector(to_unsigned( 58 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=68 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),
                    1 => std_logic_vector(to_unsigned( 121 , 8)),
                    2 => std_logic_vector(to_unsigned( 15 , 8)),
                    3 => std_logic_vector(to_unsigned( 8 , 8)),
                    4 => std_logic_vector(to_unsigned( 64 , 8)),
                    5 => std_logic_vector(to_unsigned( 34 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 96 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=69 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 8, 8)),
                    1 => std_logic_vector(to_unsigned( 35 , 8)),
                    2 => std_logic_vector(to_unsigned( 1 , 8)),
                    3 => std_logic_vector(to_unsigned( 29 , 8)),
                    4 => std_logic_vector(to_unsigned( 85 , 8)),
                    5 => std_logic_vector(to_unsigned( 47 , 8)),
                    6 => std_logic_vector(to_unsigned( 57 , 8)),
                    7 => std_logic_vector(to_unsigned( 110 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=70 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 8, 8)),
                    1 => std_logic_vector(to_unsigned( 35 , 8)),
                    2 => std_logic_vector(to_unsigned( 1 , 8)),
                    3 => std_logic_vector(to_unsigned( 29 , 8)),
                    4 => std_logic_vector(to_unsigned( 85 , 8)),
                    5 => std_logic_vector(to_unsigned( 47 , 8)),
                    6 => std_logic_vector(to_unsigned( 57 , 8)),
                    7 => std_logic_vector(to_unsigned( 110 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=71 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 104 , 8)),
                    2 => std_logic_vector(to_unsigned( 84 , 8)),
                    3 => std_logic_vector(to_unsigned( 76 , 8)),
                    4 => std_logic_vector(to_unsigned( 115 , 8)),
                    5 => std_logic_vector(to_unsigned( 2 , 8)),
                    6 => std_logic_vector(to_unsigned( 58 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=72 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),
                    1 => std_logic_vector(to_unsigned( 62 , 8)),
                    2 => std_logic_vector(to_unsigned( 94 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 43 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=73 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),
                    1 => std_logic_vector(to_unsigned( 62 , 8)),
                    2 => std_logic_vector(to_unsigned( 94 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 43 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=74 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 45, 8)),
                    1 => std_logic_vector(to_unsigned( 0 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 61 , 8)),
                    4 => std_logic_vector(to_unsigned( 103 , 8)),
                    5 => std_logic_vector(to_unsigned( 77 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 68 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=75 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 121 , 8)),
                    5 => std_logic_vector(to_unsigned( 116 , 8)),
                    6 => std_logic_vector(to_unsigned( 18 , 8)),
                    7 => std_logic_vector(to_unsigned( 70 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=76 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 121 , 8)),
                    5 => std_logic_vector(to_unsigned( 116 , 8)),
                    6 => std_logic_vector(to_unsigned( 18 , 8)),
                    7 => std_logic_vector(to_unsigned( 70 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=77 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),
                    1 => std_logic_vector(to_unsigned( 86 , 8)),
                    2 => std_logic_vector(to_unsigned( 74 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 48 , 8)),
                    5 => std_logic_vector(to_unsigned( 117 , 8)),
                    6 => std_logic_vector(to_unsigned( 28 , 8)),
                    7 => std_logic_vector(to_unsigned( 67 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=78 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 86 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 15 , 8)),
                    7 => std_logic_vector(to_unsigned( 111 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=79 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 86 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 15 , 8)),
                    7 => std_logic_vector(to_unsigned( 111 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=80 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 48 , 8)),
                    2 => std_logic_vector(to_unsigned( 22 , 8)),
                    3 => std_logic_vector(to_unsigned( 6 , 8)),
                    4 => std_logic_vector(to_unsigned( 82 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 121 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=81 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 81, 8)),
                    1 => std_logic_vector(to_unsigned( 51 , 8)),
                    2 => std_logic_vector(to_unsigned( 26 , 8)),
                    3 => std_logic_vector(to_unsigned( 5 , 8)),
                    4 => std_logic_vector(to_unsigned( 59 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=82 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 81, 8)),
                    1 => std_logic_vector(to_unsigned( 51 , 8)),
                    2 => std_logic_vector(to_unsigned( 26 , 8)),
                    3 => std_logic_vector(to_unsigned( 5 , 8)),
                    4 => std_logic_vector(to_unsigned( 59 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=83 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 88, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 26 , 8)),
                    3 => std_logic_vector(to_unsigned( 58 , 8)),
                    4 => std_logic_vector(to_unsigned( 121 , 8)),
                    5 => std_logic_vector(to_unsigned( 20 , 8)),
                    6 => std_logic_vector(to_unsigned( 49 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=84 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),
                    1 => std_logic_vector(to_unsigned( 61 , 8)),
                    2 => std_logic_vector(to_unsigned( 70 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 39 , 8)),
                    6 => std_logic_vector(to_unsigned( 94 , 8)),
                    7 => std_logic_vector(to_unsigned( 111 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=85 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),
                    1 => std_logic_vector(to_unsigned( 61 , 8)),
                    2 => std_logic_vector(to_unsigned( 70 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 39 , 8)),
                    6 => std_logic_vector(to_unsigned( 94 , 8)),
                    7 => std_logic_vector(to_unsigned( 111 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=86 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 112 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 67 , 8)),
                    5 => std_logic_vector(to_unsigned( 83 , 8)),
                    6 => std_logic_vector(to_unsigned( 35 , 8)),
                    7 => std_logic_vector(to_unsigned( 118 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=87 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 42, 8)),
                    1 => std_logic_vector(to_unsigned( 21 , 8)),
                    2 => std_logic_vector(to_unsigned( 84 , 8)),
                    3 => std_logic_vector(to_unsigned( 95 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 122 , 8)),
                    6 => std_logic_vector(to_unsigned( 16 , 8)),
                    7 => std_logic_vector(to_unsigned( 30 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=88 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 42, 8)),
                    1 => std_logic_vector(to_unsigned( 21 , 8)),
                    2 => std_logic_vector(to_unsigned( 84 , 8)),
                    3 => std_logic_vector(to_unsigned( 95 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 122 , 8)),
                    6 => std_logic_vector(to_unsigned( 16 , 8)),
                    7 => std_logic_vector(to_unsigned( 30 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=89 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),
                    1 => std_logic_vector(to_unsigned( 48 , 8)),
                    2 => std_logic_vector(to_unsigned( 3 , 8)),
                    3 => std_logic_vector(to_unsigned( 66 , 8)),
                    4 => std_logic_vector(to_unsigned( 106 , 8)),
                    5 => std_logic_vector(to_unsigned( 88 , 8)),
                    6 => std_logic_vector(to_unsigned( 80 , 8)),
                    7 => std_logic_vector(to_unsigned( 9 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=90 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 71 , 8)),
                    2 => std_logic_vector(to_unsigned( 64 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 113 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=91 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 71 , 8)),
                    2 => std_logic_vector(to_unsigned( 64 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 113 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=92 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),
                    1 => std_logic_vector(to_unsigned( 77 , 8)),
                    2 => std_logic_vector(to_unsigned( 82 , 8)),
                    3 => std_logic_vector(to_unsigned( 40 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 1 , 8)),
                    6 => std_logic_vector(to_unsigned( 45 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=93 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 115 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 124 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 105 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 71 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=94 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 115 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 124 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 105 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 71 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=95 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 2 , 8)),
                    5 => std_logic_vector(to_unsigned( 71 , 8)),
                    6 => std_logic_vector(to_unsigned( 120 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=96 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),
                    1 => std_logic_vector(to_unsigned( 58 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 26 , 8)),
                    5 => std_logic_vector(to_unsigned( 47 , 8)),
                    6 => std_logic_vector(to_unsigned( 76 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=97 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),
                    1 => std_logic_vector(to_unsigned( 58 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 26 , 8)),
                    5 => std_logic_vector(to_unsigned( 47 , 8)),
                    6 => std_logic_vector(to_unsigned( 76 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=98 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 62 , 8)),
                    3 => std_logic_vector(to_unsigned( 114 , 8)),
                    4 => std_logic_vector(to_unsigned( 17 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 83 , 8)),
                    7 => std_logic_vector(to_unsigned( 8 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=99 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 39, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 117 , 8)),
                    4 => std_logic_vector(to_unsigned( 50 , 8)),
                    5 => std_logic_vector(to_unsigned( 74 , 8)),
                    6 => std_logic_vector(to_unsigned( 91 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=100 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 39, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 117 , 8)),
                    4 => std_logic_vector(to_unsigned( 50 , 8)),
                    5 => std_logic_vector(to_unsigned( 74 , 8)),
                    6 => std_logic_vector(to_unsigned( 91 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=101 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),
                    1 => std_logic_vector(to_unsigned( 5 , 8)),
                    2 => std_logic_vector(to_unsigned( 67 , 8)),
                    3 => std_logic_vector(to_unsigned( 89 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 77 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 38 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=102 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 119 , 8)),
                    4 => std_logic_vector(to_unsigned( 104 , 8)),
                    5 => std_logic_vector(to_unsigned( 36 , 8)),
                    6 => std_logic_vector(to_unsigned( 21 , 8)),
                    7 => std_logic_vector(to_unsigned( 30 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=103 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 119 , 8)),
                    4 => std_logic_vector(to_unsigned( 104 , 8)),
                    5 => std_logic_vector(to_unsigned( 36 , 8)),
                    6 => std_logic_vector(to_unsigned( 21 , 8)),
                    7 => std_logic_vector(to_unsigned( 30 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=104 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),
                    1 => std_logic_vector(to_unsigned( 111 , 8)),
                    2 => std_logic_vector(to_unsigned( 32 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 7 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 85 , 8)),
                    7 => std_logic_vector(to_unsigned( 66 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=105 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 114 , 8)),
                    4 => std_logic_vector(to_unsigned( 34 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 79 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=106 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 114 , 8)),
                    4 => std_logic_vector(to_unsigned( 34 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 79 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=107 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 90, 8)),
                    1 => std_logic_vector(to_unsigned( 98 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 23 , 8)),
                    4 => std_logic_vector(to_unsigned( 5 , 8)),
                    5 => std_logic_vector(to_unsigned( 39 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 94 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=108 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 42, 8)),
                    1 => std_logic_vector(to_unsigned( 79 , 8)),
                    2 => std_logic_vector(to_unsigned( 112 , 8)),
                    3 => std_logic_vector(to_unsigned( 35 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 65 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=109 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 42, 8)),
                    1 => std_logic_vector(to_unsigned( 79 , 8)),
                    2 => std_logic_vector(to_unsigned( 112 , 8)),
                    3 => std_logic_vector(to_unsigned( 35 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 65 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=110 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 73, 8)),
                    1 => std_logic_vector(to_unsigned( 81 , 8)),
                    2 => std_logic_vector(to_unsigned( 2 , 8)),
                    3 => std_logic_vector(to_unsigned( 107 , 8)),
                    4 => std_logic_vector(to_unsigned( 52 , 8)),
                    5 => std_logic_vector(to_unsigned( 17 , 8)),
                    6 => std_logic_vector(to_unsigned( 41 , 8)),
                    7 => std_logic_vector(to_unsigned( 77 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=111 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 82, 8)),
                    1 => std_logic_vector(to_unsigned( 123 , 8)),
                    2 => std_logic_vector(to_unsigned( 90 , 8)),
                    3 => std_logic_vector(to_unsigned( 119 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 19 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 31 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=112 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 82, 8)),
                    1 => std_logic_vector(to_unsigned( 123 , 8)),
                    2 => std_logic_vector(to_unsigned( 90 , 8)),
                    3 => std_logic_vector(to_unsigned( 119 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 19 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 31 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=113 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 38, 8)),
                    1 => std_logic_vector(to_unsigned( 27 , 8)),
                    2 => std_logic_vector(to_unsigned( 61 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 78 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 82 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=114 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 20, 8)),
                    1 => std_logic_vector(to_unsigned( 42 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 69 , 8)),
                    4 => std_logic_vector(to_unsigned( 64 , 8)),
                    5 => std_logic_vector(to_unsigned( 60 , 8)),
                    6 => std_logic_vector(to_unsigned( 97 , 8)),
                    7 => std_logic_vector(to_unsigned( 35 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=115 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 20, 8)),
                    1 => std_logic_vector(to_unsigned( 42 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 69 , 8)),
                    4 => std_logic_vector(to_unsigned( 64 , 8)),
                    5 => std_logic_vector(to_unsigned( 60 , 8)),
                    6 => std_logic_vector(to_unsigned( 97 , 8)),
                    7 => std_logic_vector(to_unsigned( 35 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=116 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),
                    1 => std_logic_vector(to_unsigned( 96 , 8)),
                    2 => std_logic_vector(to_unsigned( 75 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 79 , 8)),
                    5 => std_logic_vector(to_unsigned( 20 , 8)),
                    6 => std_logic_vector(to_unsigned( 16 , 8)),
                    7 => std_logic_vector(to_unsigned( 69 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=117 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 101 , 8)),
                    4 => std_logic_vector(to_unsigned( 10 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 65 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=118 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 101 , 8)),
                    4 => std_logic_vector(to_unsigned( 10 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 65 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=119 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),
                    1 => std_logic_vector(to_unsigned( 7 , 8)),
                    2 => std_logic_vector(to_unsigned( 102 , 8)),
                    3 => std_logic_vector(to_unsigned( 107 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 85 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=120 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),
                    1 => std_logic_vector(to_unsigned( 99 , 8)),
                    2 => std_logic_vector(to_unsigned( 68 , 8)),
                    3 => std_logic_vector(to_unsigned( 19 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 10 , 8)),
                    6 => std_logic_vector(to_unsigned( 36 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=121 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),
                    1 => std_logic_vector(to_unsigned( 99 , 8)),
                    2 => std_logic_vector(to_unsigned( 68 , 8)),
                    3 => std_logic_vector(to_unsigned( 19 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 10 , 8)),
                    6 => std_logic_vector(to_unsigned( 36 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=122 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 81 , 8)),
                    3 => std_logic_vector(to_unsigned( 102 , 8)),
                    4 => std_logic_vector(to_unsigned( 118 , 8)),
                    5 => std_logic_vector(to_unsigned( 30 , 8)),
                    6 => std_logic_vector(to_unsigned( 63 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=123 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 19 , 8)),
                    4 => std_logic_vector(to_unsigned( 83 , 8)),
                    5 => std_logic_vector(to_unsigned( 48 , 8)),
                    6 => std_logic_vector(to_unsigned( 10 , 8)),
                    7 => std_logic_vector(to_unsigned( 31 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=124 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 19 , 8)),
                    4 => std_logic_vector(to_unsigned( 83 , 8)),
                    5 => std_logic_vector(to_unsigned( 48 , 8)),
                    6 => std_logic_vector(to_unsigned( 10 , 8)),
                    7 => std_logic_vector(to_unsigned( 31 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=125 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),
                    1 => std_logic_vector(to_unsigned( 32 , 8)),
                    2 => std_logic_vector(to_unsigned( 99 , 8)),
                    3 => std_logic_vector(to_unsigned( 16 , 8)),
                    4 => std_logic_vector(to_unsigned( 86 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 91 , 8)),
                    7 => std_logic_vector(to_unsigned( 105 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=126 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),
                    1 => std_logic_vector(to_unsigned( 108 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 14 , 8)),
                    4 => std_logic_vector(to_unsigned( 98 , 8)),
                    5 => std_logic_vector(to_unsigned( 45 , 8)),
                    6 => std_logic_vector(to_unsigned( 25 , 8)),
                    7 => std_logic_vector(to_unsigned( 35 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=127 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),
                    1 => std_logic_vector(to_unsigned( 108 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 14 , 8)),
                    4 => std_logic_vector(to_unsigned( 98 , 8)),
                    5 => std_logic_vector(to_unsigned( 45 , 8)),
                    6 => std_logic_vector(to_unsigned( 25 , 8)),
                    7 => std_logic_vector(to_unsigned( 35 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=128 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 84, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 29 , 8)),
                    3 => std_logic_vector(to_unsigned( 63 , 8)),
                    4 => std_logic_vector(to_unsigned( 45 , 8)),
                    5 => std_logic_vector(to_unsigned( 25 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 17 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=129 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 33, 8)),
                    1 => std_logic_vector(to_unsigned( 46 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 77 , 8)),
                    4 => std_logic_vector(to_unsigned( 11 , 8)),
                    5 => std_logic_vector(to_unsigned( 103 , 8)),
                    6 => std_logic_vector(to_unsigned( 116 , 8)),
                    7 => std_logic_vector(to_unsigned( 110 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=130 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 33, 8)),
                    1 => std_logic_vector(to_unsigned( 46 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 77 , 8)),
                    4 => std_logic_vector(to_unsigned( 11 , 8)),
                    5 => std_logic_vector(to_unsigned( 103 , 8)),
                    6 => std_logic_vector(to_unsigned( 116 , 8)),
                    7 => std_logic_vector(to_unsigned( 110 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=131 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 102 , 8)),
                    3 => std_logic_vector(to_unsigned( 5 , 8)),
                    4 => std_logic_vector(to_unsigned( 42 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 89 , 8)),
                    7 => std_logic_vector(to_unsigned( 77 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=132 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 15 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 80 , 8)),
                    5 => std_logic_vector(to_unsigned( 116 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 21 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=133 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 15 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 80 , 8)),
                    5 => std_logic_vector(to_unsigned( 116 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 21 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=134 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 84 , 8)),
                    3 => std_logic_vector(to_unsigned( 104 , 8)),
                    4 => std_logic_vector(to_unsigned( 54 , 8)),
                    5 => std_logic_vector(to_unsigned( 100 , 8)),
                    6 => std_logic_vector(to_unsigned( 88 , 8)),
                    7 => std_logic_vector(to_unsigned( 8 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=135 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),
                    1 => std_logic_vector(to_unsigned( 61 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 37 , 8)),
                    4 => std_logic_vector(to_unsigned( 53 , 8)),
                    5 => std_logic_vector(to_unsigned( 21 , 8)),
                    6 => std_logic_vector(to_unsigned( 114 , 8)),
                    7 => std_logic_vector(to_unsigned( 65 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=136 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),
                    1 => std_logic_vector(to_unsigned( 61 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 37 , 8)),
                    4 => std_logic_vector(to_unsigned( 53 , 8)),
                    5 => std_logic_vector(to_unsigned( 21 , 8)),
                    6 => std_logic_vector(to_unsigned( 114 , 8)),
                    7 => std_logic_vector(to_unsigned( 65 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=137 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 58, 8)),
                    1 => std_logic_vector(to_unsigned( 71 , 8)),
                    2 => std_logic_vector(to_unsigned( 43 , 8)),
                    3 => std_logic_vector(to_unsigned( 67 , 8)),
                    4 => std_logic_vector(to_unsigned( 17 , 8)),
                    5 => std_logic_vector(to_unsigned( 109 , 8)),
                    6 => std_logic_vector(to_unsigned( 80 , 8)),
                    7 => std_logic_vector(to_unsigned( 103 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=138 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 33, 8)),
                    1 => std_logic_vector(to_unsigned( 114 , 8)),
                    2 => std_logic_vector(to_unsigned( 6 , 8)),
                    3 => std_logic_vector(to_unsigned( 101 , 8)),
                    4 => std_logic_vector(to_unsigned( 55 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 45 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=139 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 33, 8)),
                    1 => std_logic_vector(to_unsigned( 114 , 8)),
                    2 => std_logic_vector(to_unsigned( 6 , 8)),
                    3 => std_logic_vector(to_unsigned( 101 , 8)),
                    4 => std_logic_vector(to_unsigned( 55 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 45 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=140 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 48 , 8)),
                    2 => std_logic_vector(to_unsigned( 59 , 8)),
                    3 => std_logic_vector(to_unsigned( 81 , 8)),
                    4 => std_logic_vector(to_unsigned( 12 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 110 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=141 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 24 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 110 , 8)),
                    5 => std_logic_vector(to_unsigned( 1 , 8)),
                    6 => std_logic_vector(to_unsigned( 5 , 8)),
                    7 => std_logic_vector(to_unsigned( 57 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=142 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 24 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 110 , 8)),
                    5 => std_logic_vector(to_unsigned( 1 , 8)),
                    6 => std_logic_vector(to_unsigned( 5 , 8)),
                    7 => std_logic_vector(to_unsigned( 57 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=143 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 40 , 8)),
                    3 => std_logic_vector(to_unsigned( 18 , 8)),
                    4 => std_logic_vector(to_unsigned( 23 , 8)),
                    5 => std_logic_vector(to_unsigned( 35 , 8)),
                    6 => std_logic_vector(to_unsigned( 30 , 8)),
                    7 => std_logic_vector(to_unsigned( 113 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=144 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 51 , 8)),
                    2 => std_logic_vector(to_unsigned( 114 , 8)),
                    3 => std_logic_vector(to_unsigned( 67 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 62 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=145 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 51 , 8)),
                    2 => std_logic_vector(to_unsigned( 114 , 8)),
                    3 => std_logic_vector(to_unsigned( 67 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 62 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=146 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 77 , 8)),
                    2 => std_logic_vector(to_unsigned( 49 , 8)),
                    3 => std_logic_vector(to_unsigned( 21 , 8)),
                    4 => std_logic_vector(to_unsigned( 17 , 8)),
                    5 => std_logic_vector(to_unsigned( 36 , 8)),
                    6 => std_logic_vector(to_unsigned( 56 , 8)),
                    7 => std_logic_vector(to_unsigned( 31 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=147 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),
                    1 => std_logic_vector(to_unsigned( 96 , 8)),
                    2 => std_logic_vector(to_unsigned( 19 , 8)),
                    3 => std_logic_vector(to_unsigned( 12 , 8)),
                    4 => std_logic_vector(to_unsigned( 26 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 7 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=148 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),
                    1 => std_logic_vector(to_unsigned( 96 , 8)),
                    2 => std_logic_vector(to_unsigned( 19 , 8)),
                    3 => std_logic_vector(to_unsigned( 12 , 8)),
                    4 => std_logic_vector(to_unsigned( 26 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 7 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=149 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 45, 8)),
                    1 => std_logic_vector(to_unsigned( 81 , 8)),
                    2 => std_logic_vector(to_unsigned( 26 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 5 , 8)),
                    5 => std_logic_vector(to_unsigned( 21 , 8)),
                    6 => std_logic_vector(to_unsigned( 76 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=150 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),
                    1 => std_logic_vector(to_unsigned( 12 , 8)),
                    2 => std_logic_vector(to_unsigned( 114 , 8)),
                    3 => std_logic_vector(to_unsigned( 93 , 8)),
                    4 => std_logic_vector(to_unsigned( 19 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=151 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),
                    1 => std_logic_vector(to_unsigned( 12 , 8)),
                    2 => std_logic_vector(to_unsigned( 114 , 8)),
                    3 => std_logic_vector(to_unsigned( 93 , 8)),
                    4 => std_logic_vector(to_unsigned( 19 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=152 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 14 , 8)),
                    2 => std_logic_vector(to_unsigned( 112 , 8)),
                    3 => std_logic_vector(to_unsigned( 21 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 82 , 8)),
                    6 => std_logic_vector(to_unsigned( 122 , 8)),
                    7 => std_logic_vector(to_unsigned( 4 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=153 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 115, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 9 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 25 , 8)),
                    5 => std_logic_vector(to_unsigned( 94 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 78 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=154 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 115, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 9 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 25 , 8)),
                    5 => std_logic_vector(to_unsigned( 94 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 78 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=155 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 63 , 8)),
                    3 => std_logic_vector(to_unsigned( 59 , 8)),
                    4 => std_logic_vector(to_unsigned( 75 , 8)),
                    5 => std_logic_vector(to_unsigned( 5 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 45 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=156 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 92 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 82 , 8)),
                    4 => std_logic_vector(to_unsigned( 10 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 27 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=157 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 92 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 82 , 8)),
                    4 => std_logic_vector(to_unsigned( 10 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 27 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=158 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),
                    1 => std_logic_vector(to_unsigned( 115 , 8)),
                    2 => std_logic_vector(to_unsigned( 52 , 8)),
                    3 => std_logic_vector(to_unsigned( 60 , 8)),
                    4 => std_logic_vector(to_unsigned( 88 , 8)),
                    5 => std_logic_vector(to_unsigned( 72 , 8)),
                    6 => std_logic_vector(to_unsigned( 94 , 8)),
                    7 => std_logic_vector(to_unsigned( 20 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=159 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 115, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 61 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 122 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 78 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=160 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 115, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 61 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 122 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 78 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=161 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 36 , 8)),
                    4 => std_logic_vector(to_unsigned( 108 , 8)),
                    5 => std_logic_vector(to_unsigned( 50 , 8)),
                    6 => std_logic_vector(to_unsigned( 28 , 8)),
                    7 => std_logic_vector(to_unsigned( 61 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=162 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 110 , 8)),
                    2 => std_logic_vector(to_unsigned( 57 , 8)),
                    3 => std_logic_vector(to_unsigned( 27 , 8)),
                    4 => std_logic_vector(to_unsigned( 65 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 23 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=163 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 110 , 8)),
                    2 => std_logic_vector(to_unsigned( 57 , 8)),
                    3 => std_logic_vector(to_unsigned( 27 , 8)),
                    4 => std_logic_vector(to_unsigned( 65 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 23 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=164 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 115, 8)),
                    1 => std_logic_vector(to_unsigned( 59 , 8)),
                    2 => std_logic_vector(to_unsigned( 100 , 8)),
                    3 => std_logic_vector(to_unsigned( 106 , 8)),
                    4 => std_logic_vector(to_unsigned( 54 , 8)),
                    5 => std_logic_vector(to_unsigned( 42 , 8)),
                    6 => std_logic_vector(to_unsigned( 10 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=165 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),
                    1 => std_logic_vector(to_unsigned( 99 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 113 , 8)),
                    4 => std_logic_vector(to_unsigned( 63 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 12 , 8)),
                    7 => std_logic_vector(to_unsigned( 45 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=166 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),
                    1 => std_logic_vector(to_unsigned( 99 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 113 , 8)),
                    4 => std_logic_vector(to_unsigned( 63 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 12 , 8)),
                    7 => std_logic_vector(to_unsigned( 45 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=167 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 105 , 8)),
                    2 => std_logic_vector(to_unsigned( 21 , 8)),
                    3 => std_logic_vector(to_unsigned( 114 , 8)),
                    4 => std_logic_vector(to_unsigned( 34 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 65 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=168 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 88, 8)),
                    1 => std_logic_vector(to_unsigned( 103 , 8)),
                    2 => std_logic_vector(to_unsigned( 43 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 48 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 31 , 8)),
                    7 => std_logic_vector(to_unsigned( 117 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=169 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 88, 8)),
                    1 => std_logic_vector(to_unsigned( 103 , 8)),
                    2 => std_logic_vector(to_unsigned( 43 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 48 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 31 , 8)),
                    7 => std_logic_vector(to_unsigned( 117 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=170 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 34 , 8)),
                    3 => std_logic_vector(to_unsigned( 63 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 5 , 8)),
                    6 => std_logic_vector(to_unsigned( 26 , 8)),
                    7 => std_logic_vector(to_unsigned( 100 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=171 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 106 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 51 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=172 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 106 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 51 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=173 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 63, 8)),
                    1 => std_logic_vector(to_unsigned( 52 , 8)),
                    2 => std_logic_vector(to_unsigned( 1 , 8)),
                    3 => std_logic_vector(to_unsigned( 81 , 8)),
                    4 => std_logic_vector(to_unsigned( 99 , 8)),
                    5 => std_logic_vector(to_unsigned( 15 , 8)),
                    6 => std_logic_vector(to_unsigned( 44 , 8)),
                    7 => std_logic_vector(to_unsigned( 70 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=174 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 62 , 8)),
                    4 => std_logic_vector(to_unsigned( 119 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 32 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=175 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 62 , 8)),
                    4 => std_logic_vector(to_unsigned( 119 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 32 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=176 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),
                    1 => std_logic_vector(to_unsigned( 104 , 8)),
                    2 => std_logic_vector(to_unsigned( 64 , 8)),
                    3 => std_logic_vector(to_unsigned( 45 , 8)),
                    4 => std_logic_vector(to_unsigned( 51 , 8)),
                    5 => std_logic_vector(to_unsigned( 83 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 98 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=177 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 77 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 34 , 8)),
                    6 => std_logic_vector(to_unsigned( 57 , 8)),
                    7 => std_logic_vector(to_unsigned( 5 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=178 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 77 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 34 , 8)),
                    6 => std_logic_vector(to_unsigned( 57 , 8)),
                    7 => std_logic_vector(to_unsigned( 5 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=179 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 105, 8)),
                    1 => std_logic_vector(to_unsigned( 23 , 8)),
                    2 => std_logic_vector(to_unsigned( 61 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 72 , 8)),
                    5 => std_logic_vector(to_unsigned( 36 , 8)),
                    6 => std_logic_vector(to_unsigned( 66 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=180 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 74 , 8)),
                    3 => std_logic_vector(to_unsigned( 122 , 8)),
                    4 => std_logic_vector(to_unsigned( 104 , 8)),
                    5 => std_logic_vector(to_unsigned( 56 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=181 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 74 , 8)),
                    3 => std_logic_vector(to_unsigned( 122 , 8)),
                    4 => std_logic_vector(to_unsigned( 104 , 8)),
                    5 => std_logic_vector(to_unsigned( 56 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=182 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),
                    1 => std_logic_vector(to_unsigned( 17 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 84 , 8)),
                    4 => std_logic_vector(to_unsigned( 22 , 8)),
                    5 => std_logic_vector(to_unsigned( 55 , 8)),
                    6 => std_logic_vector(to_unsigned( 97 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=183 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 101 , 8)),
                    3 => std_logic_vector(to_unsigned( 21 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 41 , 8)),
                    6 => std_logic_vector(to_unsigned( 7 , 8)),
                    7 => std_logic_vector(to_unsigned( 96 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=184 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 101 , 8)),
                    3 => std_logic_vector(to_unsigned( 21 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 41 , 8)),
                    6 => std_logic_vector(to_unsigned( 7 , 8)),
                    7 => std_logic_vector(to_unsigned( 96 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=185 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 117 , 8)),
                    2 => std_logic_vector(to_unsigned( 83 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 5 , 8)),
                    5 => std_logic_vector(to_unsigned( 12 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 97 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=186 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 16, 8)),
                    1 => std_logic_vector(to_unsigned( 93 , 8)),
                    2 => std_logic_vector(to_unsigned( 28 , 8)),
                    3 => std_logic_vector(to_unsigned( 114 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 81 , 8)),
                    7 => std_logic_vector(to_unsigned( 101 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=187 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 16, 8)),
                    1 => std_logic_vector(to_unsigned( 93 , 8)),
                    2 => std_logic_vector(to_unsigned( 28 , 8)),
                    3 => std_logic_vector(to_unsigned( 114 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 81 , 8)),
                    7 => std_logic_vector(to_unsigned( 101 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=188 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 118, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 53 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 87 , 8)),
                    6 => std_logic_vector(to_unsigned( 114 , 8)),
                    7 => std_logic_vector(to_unsigned( 71 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=189 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 5 , 8)),
                    2 => std_logic_vector(to_unsigned( 39 , 8)),
                    3 => std_logic_vector(to_unsigned( 20 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 15 , 8)),
                    6 => std_logic_vector(to_unsigned( 82 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=190 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 5 , 8)),
                    2 => std_logic_vector(to_unsigned( 39 , 8)),
                    3 => std_logic_vector(to_unsigned( 20 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 15 , 8)),
                    6 => std_logic_vector(to_unsigned( 82 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=191 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),
                    1 => std_logic_vector(to_unsigned( 58 , 8)),
                    2 => std_logic_vector(to_unsigned( 36 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 99 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 122 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=192 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 113, 8)),
                    1 => std_logic_vector(to_unsigned( 59 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 55 , 8)),
                    4 => std_logic_vector(to_unsigned( 50 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 117 , 8)),
                    7 => std_logic_vector(to_unsigned( 30 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=193 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 113, 8)),
                    1 => std_logic_vector(to_unsigned( 59 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 55 , 8)),
                    4 => std_logic_vector(to_unsigned( 50 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 117 , 8)),
                    7 => std_logic_vector(to_unsigned( 30 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=194 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 47, 8)),
                    1 => std_logic_vector(to_unsigned( 119 , 8)),
                    2 => std_logic_vector(to_unsigned( 57 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 65 , 8)),
                    5 => std_logic_vector(to_unsigned( 103 , 8)),
                    6 => std_logic_vector(to_unsigned( 35 , 8)),
                    7 => std_logic_vector(to_unsigned( 69 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=195 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 41, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 75 , 8)),
                    3 => std_logic_vector(to_unsigned( 92 , 8)),
                    4 => std_logic_vector(to_unsigned( 86 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 64 , 8)),
                    7 => std_logic_vector(to_unsigned( 56 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=196 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 41, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 75 , 8)),
                    3 => std_logic_vector(to_unsigned( 92 , 8)),
                    4 => std_logic_vector(to_unsigned( 86 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 64 , 8)),
                    7 => std_logic_vector(to_unsigned( 56 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=197 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),
                    1 => std_logic_vector(to_unsigned( 45 , 8)),
                    2 => std_logic_vector(to_unsigned( 64 , 8)),
                    3 => std_logic_vector(to_unsigned( 73 , 8)),
                    4 => std_logic_vector(to_unsigned( 87 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=198 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 109, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 2 , 8)),
                    3 => std_logic_vector(to_unsigned( 115 , 8)),
                    4 => std_logic_vector(to_unsigned( 42 , 8)),
                    5 => std_logic_vector(to_unsigned( 37 , 8)),
                    6 => std_logic_vector(to_unsigned( 105 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=199 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 109, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 2 , 8)),
                    3 => std_logic_vector(to_unsigned( 115 , 8)),
                    4 => std_logic_vector(to_unsigned( 42 , 8)),
                    5 => std_logic_vector(to_unsigned( 37 , 8)),
                    6 => std_logic_vector(to_unsigned( 105 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=200 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 73, 8)),
                    1 => std_logic_vector(to_unsigned( 44 , 8)),
                    2 => std_logic_vector(to_unsigned( 94 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 20 , 8)),
                    6 => std_logic_vector(to_unsigned( 116 , 8)),
                    7 => std_logic_vector(to_unsigned( 120 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=201 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 33 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 28 , 8)),
                    4 => std_logic_vector(to_unsigned( 68 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 94 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=202 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 33 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 28 , 8)),
                    4 => std_logic_vector(to_unsigned( 68 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 94 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=203 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 89 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 31 , 8)),
                    4 => std_logic_vector(to_unsigned( 41 , 8)),
                    5 => std_logic_vector(to_unsigned( 74 , 8)),
                    6 => std_logic_vector(to_unsigned( 79 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=204 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 68 , 8)),
                    2 => std_logic_vector(to_unsigned( 51 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 5 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 56 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=205 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 68 , 8)),
                    2 => std_logic_vector(to_unsigned( 51 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 5 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 56 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=206 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 104 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 27 , 8)),
                    5 => std_logic_vector(to_unsigned( 15 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=207 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 26 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 52 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=208 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 26 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 52 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=209 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 19 , 8)),
                    2 => std_logic_vector(to_unsigned( 79 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 41 , 8)),
                    5 => std_logic_vector(to_unsigned( 7 , 8)),
                    6 => std_logic_vector(to_unsigned( 89 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=210 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 11 , 8)),
                    3 => std_logic_vector(to_unsigned( 109 , 8)),
                    4 => std_logic_vector(to_unsigned( 84 , 8)),
                    5 => std_logic_vector(to_unsigned( 117 , 8)),
                    6 => std_logic_vector(to_unsigned( 44 , 8)),
                    7 => std_logic_vector(to_unsigned( 122 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=211 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 11 , 8)),
                    3 => std_logic_vector(to_unsigned( 109 , 8)),
                    4 => std_logic_vector(to_unsigned( 84 , 8)),
                    5 => std_logic_vector(to_unsigned( 117 , 8)),
                    6 => std_logic_vector(to_unsigned( 44 , 8)),
                    7 => std_logic_vector(to_unsigned( 122 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=212 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 12, 8)),
                    1 => std_logic_vector(to_unsigned( 86 , 8)),
                    2 => std_logic_vector(to_unsigned( 30 , 8)),
                    3 => std_logic_vector(to_unsigned( 103 , 8)),
                    4 => std_logic_vector(to_unsigned( 40 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 49 , 8)),
                    7 => std_logic_vector(to_unsigned( 19 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=213 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=214 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=215 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 51, 8)),
                    1 => std_logic_vector(to_unsigned( 96 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 67 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 29 , 8)),
                    7 => std_logic_vector(to_unsigned( 13 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=216 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),
                    1 => std_logic_vector(to_unsigned( 45 , 8)),
                    2 => std_logic_vector(to_unsigned( 83 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 72 , 8)),
                    5 => std_logic_vector(to_unsigned( 64 , 8)),
                    6 => std_logic_vector(to_unsigned( 35 , 8)),
                    7 => std_logic_vector(to_unsigned( 122 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=217 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),
                    1 => std_logic_vector(to_unsigned( 45 , 8)),
                    2 => std_logic_vector(to_unsigned( 83 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 72 , 8)),
                    5 => std_logic_vector(to_unsigned( 64 , 8)),
                    6 => std_logic_vector(to_unsigned( 35 , 8)),
                    7 => std_logic_vector(to_unsigned( 122 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=218 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 101 , 8)),
                    2 => std_logic_vector(to_unsigned( 81 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 97 , 8)),
                    5 => std_logic_vector(to_unsigned( 71 , 8)),
                    6 => std_logic_vector(to_unsigned( 61 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=219 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 53 , 8)),
                    3 => std_logic_vector(to_unsigned( 99 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 5 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 115 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=220 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 53 , 8)),
                    3 => std_logic_vector(to_unsigned( 99 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 5 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 115 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=221 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),
                    1 => std_logic_vector(to_unsigned( 45 , 8)),
                    2 => std_logic_vector(to_unsigned( 90 , 8)),
                    3 => std_logic_vector(to_unsigned( 65 , 8)),
                    4 => std_logic_vector(to_unsigned( 40 , 8)),
                    5 => std_logic_vector(to_unsigned( 0 , 8)),
                    6 => std_logic_vector(to_unsigned( 72 , 8)),
                    7 => std_logic_vector(to_unsigned( 113 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=222 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 57 , 8)),
                    2 => std_logic_vector(to_unsigned( 21 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 94 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=223 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 57 , 8)),
                    2 => std_logic_vector(to_unsigned( 21 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 94 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=224 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 99, 8)),
                    1 => std_logic_vector(to_unsigned( 86 , 8)),
                    2 => std_logic_vector(to_unsigned( 74 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 28 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 122 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=225 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 76, 8)),
                    1 => std_logic_vector(to_unsigned( 17 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 29 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 70 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=226 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 76, 8)),
                    1 => std_logic_vector(to_unsigned( 17 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 29 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 70 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=227 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 101 , 8)),
                    2 => std_logic_vector(to_unsigned( 56 , 8)),
                    3 => std_logic_vector(to_unsigned( 28 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 119 , 8)),
                    6 => std_logic_vector(to_unsigned( 80 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=228 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 33 , 8)),
                    2 => std_logic_vector(to_unsigned( 69 , 8)),
                    3 => std_logic_vector(to_unsigned( 53 , 8)),
                    4 => std_logic_vector(to_unsigned( 9 , 8)),
                    5 => std_logic_vector(to_unsigned( 124 , 8)),
                    6 => std_logic_vector(to_unsigned( 94 , 8)),
                    7 => std_logic_vector(to_unsigned( 25 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=229 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 33 , 8)),
                    2 => std_logic_vector(to_unsigned( 69 , 8)),
                    3 => std_logic_vector(to_unsigned( 53 , 8)),
                    4 => std_logic_vector(to_unsigned( 9 , 8)),
                    5 => std_logic_vector(to_unsigned( 124 , 8)),
                    6 => std_logic_vector(to_unsigned( 94 , 8)),
                    7 => std_logic_vector(to_unsigned( 25 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=230 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 38, 8)),
                    1 => std_logic_vector(to_unsigned( 81 , 8)),
                    2 => std_logic_vector(to_unsigned( 112 , 8)),
                    3 => std_logic_vector(to_unsigned( 43 , 8)),
                    4 => std_logic_vector(to_unsigned( 23 , 8)),
                    5 => std_logic_vector(to_unsigned( 105 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 70 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=231 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),
                    1 => std_logic_vector(to_unsigned( 32 , 8)),
                    2 => std_logic_vector(to_unsigned( 65 , 8)),
                    3 => std_logic_vector(to_unsigned( 122 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 84 , 8)),
                    6 => std_logic_vector(to_unsigned( 79 , 8)),
                    7 => std_logic_vector(to_unsigned( 1 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=232 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),
                    1 => std_logic_vector(to_unsigned( 32 , 8)),
                    2 => std_logic_vector(to_unsigned( 65 , 8)),
                    3 => std_logic_vector(to_unsigned( 122 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 84 , 8)),
                    6 => std_logic_vector(to_unsigned( 79 , 8)),
                    7 => std_logic_vector(to_unsigned( 1 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=233 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 54, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 31 , 8)),
                    3 => std_logic_vector(to_unsigned( 18 , 8)),
                    4 => std_logic_vector(to_unsigned( 79 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 73 , 8)),
                    7 => std_logic_vector(to_unsigned( 120 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=234 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 45 , 8)),
                    3 => std_logic_vector(to_unsigned( 16 , 8)),
                    4 => std_logic_vector(to_unsigned( 94 , 8)),
                    5 => std_logic_vector(to_unsigned( 33 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 12 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=235 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 45 , 8)),
                    3 => std_logic_vector(to_unsigned( 16 , 8)),
                    4 => std_logic_vector(to_unsigned( 94 , 8)),
                    5 => std_logic_vector(to_unsigned( 33 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 12 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=236 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 3 , 8)),
                    2 => std_logic_vector(to_unsigned( 103 , 8)),
                    3 => std_logic_vector(to_unsigned( 86 , 8)),
                    4 => std_logic_vector(to_unsigned( 79 , 8)),
                    5 => std_logic_vector(to_unsigned( 64 , 8)),
                    6 => std_logic_vector(to_unsigned( 91 , 8)),
                    7 => std_logic_vector(to_unsigned( 68 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=237 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),
                    1 => std_logic_vector(to_unsigned( 68 , 8)),
                    2 => std_logic_vector(to_unsigned( 30 , 8)),
                    3 => std_logic_vector(to_unsigned( 91 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 41 , 8)),
                    6 => std_logic_vector(to_unsigned( 113 , 8)),
                    7 => std_logic_vector(to_unsigned( 75 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=238 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),
                    1 => std_logic_vector(to_unsigned( 68 , 8)),
                    2 => std_logic_vector(to_unsigned( 30 , 8)),
                    3 => std_logic_vector(to_unsigned( 91 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 41 , 8)),
                    6 => std_logic_vector(to_unsigned( 113 , 8)),
                    7 => std_logic_vector(to_unsigned( 75 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=239 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),
                    1 => std_logic_vector(to_unsigned( 35 , 8)),
                    2 => std_logic_vector(to_unsigned( 43 , 8)),
                    3 => std_logic_vector(to_unsigned( 25 , 8)),
                    4 => std_logic_vector(to_unsigned( 53 , 8)),
                    5 => std_logic_vector(to_unsigned( 13 , 8)),
                    6 => std_logic_vector(to_unsigned( 19 , 8)),
                    7 => std_logic_vector(to_unsigned( 122 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=240 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 72, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 105 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 53 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=241 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 72, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 105 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 53 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=242 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 35 , 8)),
                    2 => std_logic_vector(to_unsigned( 65 , 8)),
                    3 => std_logic_vector(to_unsigned( 17 , 8)),
                    4 => std_logic_vector(to_unsigned( 105 , 8)),
                    5 => std_logic_vector(to_unsigned( 77 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=243 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),
                    1 => std_logic_vector(to_unsigned( 90 , 8)),
                    2 => std_logic_vector(to_unsigned( 105 , 8)),
                    3 => std_logic_vector(to_unsigned( 36 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 77 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=244 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),
                    1 => std_logic_vector(to_unsigned( 90 , 8)),
                    2 => std_logic_vector(to_unsigned( 105 , 8)),
                    3 => std_logic_vector(to_unsigned( 36 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 77 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=245 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),
                    1 => std_logic_vector(to_unsigned( 40 , 8)),
                    2 => std_logic_vector(to_unsigned( 13 , 8)),
                    3 => std_logic_vector(to_unsigned( 104 , 8)),
                    4 => std_logic_vector(to_unsigned( 3 , 8)),
                    5 => std_logic_vector(to_unsigned( 121 , 8)),
                    6 => std_logic_vector(to_unsigned( 50 , 8)),
                    7 => std_logic_vector(to_unsigned( 88 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=246 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),
                    1 => std_logic_vector(to_unsigned( 91 , 8)),
                    2 => std_logic_vector(to_unsigned( 49 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 75 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 16 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=247 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),
                    1 => std_logic_vector(to_unsigned( 91 , 8)),
                    2 => std_logic_vector(to_unsigned( 49 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 75 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 16 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=248 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 77, 8)),
                    1 => std_logic_vector(to_unsigned( 124 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 56 , 8)),
                    4 => std_logic_vector(to_unsigned( 103 , 8)),
                    5 => std_logic_vector(to_unsigned( 119 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 21 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=249 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 49 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 102 , 8)),
                    7 => std_logic_vector(to_unsigned( 42 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=250 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 49 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 102 , 8)),
                    7 => std_logic_vector(to_unsigned( 42 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=251 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),
                    1 => std_logic_vector(to_unsigned( 79 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 99 , 8)),
                    4 => std_logic_vector(to_unsigned( 2 , 8)),
                    5 => std_logic_vector(to_unsigned( 112 , 8)),
                    6 => std_logic_vector(to_unsigned( 67 , 8)),
                    7 => std_logic_vector(to_unsigned( 117 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=252 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 46 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 66 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 80 , 8)),
                    7 => std_logic_vector(to_unsigned( 74 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=253 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 46 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 66 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 80 , 8)),
                    7 => std_logic_vector(to_unsigned( 74 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=254 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 8, 8)),
                    1 => std_logic_vector(to_unsigned( 98 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 14 , 8)),
                    4 => std_logic_vector(to_unsigned( 34 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 78 , 8)),
                    7 => std_logic_vector(to_unsigned( 45 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=255 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 76, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 66 , 8)),
                    4 => std_logic_vector(to_unsigned( 34 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 88 , 8)),
                    7 => std_logic_vector(to_unsigned( 1 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=256 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 76, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 66 , 8)),
                    4 => std_logic_vector(to_unsigned( 34 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 88 , 8)),
                    7 => std_logic_vector(to_unsigned( 1 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=257 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),
                    1 => std_logic_vector(to_unsigned( 100 , 8)),
                    2 => std_logic_vector(to_unsigned( 35 , 8)),
                    3 => std_logic_vector(to_unsigned( 112 , 8)),
                    4 => std_logic_vector(to_unsigned( 73 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 87 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=258 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 84, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 8 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 64 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=259 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 84, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 8 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 64 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=260 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 51 , 8)),
                    3 => std_logic_vector(to_unsigned( 45 , 8)),
                    4 => std_logic_vector(to_unsigned( 123 , 8)),
                    5 => std_logic_vector(to_unsigned( 13 , 8)),
                    6 => std_logic_vector(to_unsigned( 57 , 8)),
                    7 => std_logic_vector(to_unsigned( 87 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=261 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 121 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 39 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 0 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=262 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 121 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 39 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 0 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=263 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 103 , 8)),
                    2 => std_logic_vector(to_unsigned( 90 , 8)),
                    3 => std_logic_vector(to_unsigned( 37 , 8)),
                    4 => std_logic_vector(to_unsigned( 19 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 54 , 8)),
                    7 => std_logic_vector(to_unsigned( 15 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=264 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 103 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 12 , 8)),
                    5 => std_logic_vector(to_unsigned( 95 , 8)),
                    6 => std_logic_vector(to_unsigned( 67 , 8)),
                    7 => std_logic_vector(to_unsigned( 113 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=265 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 103 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 12 , 8)),
                    5 => std_logic_vector(to_unsigned( 95 , 8)),
                    6 => std_logic_vector(to_unsigned( 67 , 8)),
                    7 => std_logic_vector(to_unsigned( 113 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=266 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 17, 8)),
                    1 => std_logic_vector(to_unsigned( 123 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 99 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 84 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 23 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=267 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 30 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 21 , 8)),
                    7 => std_logic_vector(to_unsigned( 101 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=268 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 30 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 21 , 8)),
                    7 => std_logic_vector(to_unsigned( 101 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=269 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 12, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 23 , 8)),
                    3 => std_logic_vector(to_unsigned( 111 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 42 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=270 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 97, 8)),
                    1 => std_logic_vector(to_unsigned( 92 , 8)),
                    2 => std_logic_vector(to_unsigned( 34 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 53 , 8)),
                    5 => std_logic_vector(to_unsigned( 45 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 81 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=271 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 97, 8)),
                    1 => std_logic_vector(to_unsigned( 92 , 8)),
                    2 => std_logic_vector(to_unsigned( 34 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 53 , 8)),
                    5 => std_logic_vector(to_unsigned( 45 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 81 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=272 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),
                    1 => std_logic_vector(to_unsigned( 39 , 8)),
                    2 => std_logic_vector(to_unsigned( 56 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 68 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 74 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=273 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 118 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 38 , 8)),
                    5 => std_logic_vector(to_unsigned( 109 , 8)),
                    6 => std_logic_vector(to_unsigned( 32 , 8)),
                    7 => std_logic_vector(to_unsigned( 96 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=274 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 118 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 38 , 8)),
                    5 => std_logic_vector(to_unsigned( 109 , 8)),
                    6 => std_logic_vector(to_unsigned( 32 , 8)),
                    7 => std_logic_vector(to_unsigned( 96 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=275 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 46, 8)),
                    1 => std_logic_vector(to_unsigned( 18 , 8)),
                    2 => std_logic_vector(to_unsigned( 71 , 8)),
                    3 => std_logic_vector(to_unsigned( 111 , 8)),
                    4 => std_logic_vector(to_unsigned( 26 , 8)),
                    5 => std_logic_vector(to_unsigned( 84 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=276 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),
                    1 => std_logic_vector(to_unsigned( 66 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 56 , 8)),
                    5 => std_logic_vector(to_unsigned( 62 , 8)),
                    6 => std_logic_vector(to_unsigned( 13 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=277 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),
                    1 => std_logic_vector(to_unsigned( 66 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 56 , 8)),
                    5 => std_logic_vector(to_unsigned( 62 , 8)),
                    6 => std_logic_vector(to_unsigned( 13 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=278 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 89 , 8)),
                    2 => std_logic_vector(to_unsigned( 85 , 8)),
                    3 => std_logic_vector(to_unsigned( 117 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 21 , 8)),
                    6 => std_logic_vector(to_unsigned( 52 , 8)),
                    7 => std_logic_vector(to_unsigned( 36 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=279 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 46, 8)),
                    1 => std_logic_vector(to_unsigned( 42 , 8)),
                    2 => std_logic_vector(to_unsigned( 117 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 124 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=280 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 46, 8)),
                    1 => std_logic_vector(to_unsigned( 42 , 8)),
                    2 => std_logic_vector(to_unsigned( 117 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 124 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=281 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 118, 8)),
                    1 => std_logic_vector(to_unsigned( 34 , 8)),
                    2 => std_logic_vector(to_unsigned( 64 , 8)),
                    3 => std_logic_vector(to_unsigned( 103 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 76 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 88 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=282 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 46 , 8)),
                    2 => std_logic_vector(to_unsigned( 18 , 8)),
                    3 => std_logic_vector(to_unsigned( 53 , 8)),
                    4 => std_logic_vector(to_unsigned( 37 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=283 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 46 , 8)),
                    2 => std_logic_vector(to_unsigned( 18 , 8)),
                    3 => std_logic_vector(to_unsigned( 53 , 8)),
                    4 => std_logic_vector(to_unsigned( 37 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=284 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),
                    1 => std_logic_vector(to_unsigned( 62 , 8)),
                    2 => std_logic_vector(to_unsigned( 27 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 78 , 8)),
                    5 => std_logic_vector(to_unsigned( 35 , 8)),
                    6 => std_logic_vector(to_unsigned( 105 , 8)),
                    7 => std_logic_vector(to_unsigned( 94 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=285 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 34 , 8)),
                    2 => std_logic_vector(to_unsigned( 81 , 8)),
                    3 => std_logic_vector(to_unsigned( 66 , 8)),
                    4 => std_logic_vector(to_unsigned( 76 , 8)),
                    5 => std_logic_vector(to_unsigned( 30 , 8)),
                    6 => std_logic_vector(to_unsigned( 41 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=286 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 34 , 8)),
                    2 => std_logic_vector(to_unsigned( 81 , 8)),
                    3 => std_logic_vector(to_unsigned( 66 , 8)),
                    4 => std_logic_vector(to_unsigned( 76 , 8)),
                    5 => std_logic_vector(to_unsigned( 30 , 8)),
                    6 => std_logic_vector(to_unsigned( 41 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=287 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),
                    1 => std_logic_vector(to_unsigned( 12 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 70 , 8)),
                    4 => std_logic_vector(to_unsigned( 32 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 23 , 8)),
                    7 => std_logic_vector(to_unsigned( 36 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=288 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 32 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 25 , 8)),
                    5 => std_logic_vector(to_unsigned( 19 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 58 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=289 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 32 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 25 , 8)),
                    5 => std_logic_vector(to_unsigned( 19 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 58 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=290 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 106, 8)),
                    1 => std_logic_vector(to_unsigned( 119 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 84 , 8)),
                    4 => std_logic_vector(to_unsigned( 123 , 8)),
                    5 => std_logic_vector(to_unsigned( 48 , 8)),
                    6 => std_logic_vector(to_unsigned( 77 , 8)),
                    7 => std_logic_vector(to_unsigned( 13 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=291 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),
                    1 => std_logic_vector(to_unsigned( 54 , 8)),
                    2 => std_logic_vector(to_unsigned( 46 , 8)),
                    3 => std_logic_vector(to_unsigned( 96 , 8)),
                    4 => std_logic_vector(to_unsigned( 64 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=292 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),
                    1 => std_logic_vector(to_unsigned( 54 , 8)),
                    2 => std_logic_vector(to_unsigned( 46 , 8)),
                    3 => std_logic_vector(to_unsigned( 96 , 8)),
                    4 => std_logic_vector(to_unsigned( 64 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=293 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),
                    1 => std_logic_vector(to_unsigned( 32 , 8)),
                    2 => std_logic_vector(to_unsigned( 106 , 8)),
                    3 => std_logic_vector(to_unsigned( 63 , 8)),
                    4 => std_logic_vector(to_unsigned( 88 , 8)),
                    5 => std_logic_vector(to_unsigned( 21 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 98 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=294 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 40, 8)),
                    1 => std_logic_vector(to_unsigned( 10 , 8)),
                    2 => std_logic_vector(to_unsigned( 54 , 8)),
                    3 => std_logic_vector(to_unsigned( 62 , 8)),
                    4 => std_logic_vector(to_unsigned( 21 , 8)),
                    5 => std_logic_vector(to_unsigned( 115 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 79 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=295 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 40, 8)),
                    1 => std_logic_vector(to_unsigned( 10 , 8)),
                    2 => std_logic_vector(to_unsigned( 54 , 8)),
                    3 => std_logic_vector(to_unsigned( 62 , 8)),
                    4 => std_logic_vector(to_unsigned( 21 , 8)),
                    5 => std_logic_vector(to_unsigned( 115 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 79 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=296 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 10 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 101 , 8)),
                    4 => std_logic_vector(to_unsigned( 50 , 8)),
                    5 => std_logic_vector(to_unsigned( 39 , 8)),
                    6 => std_logic_vector(to_unsigned( 23 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=297 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 103 , 8)),
                    2 => std_logic_vector(to_unsigned( 81 , 8)),
                    3 => std_logic_vector(to_unsigned( 91 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 123 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=298 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 103 , 8)),
                    2 => std_logic_vector(to_unsigned( 81 , 8)),
                    3 => std_logic_vector(to_unsigned( 91 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 123 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=299 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 56 , 8)),
                    3 => std_logic_vector(to_unsigned( 41 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 110 , 8)),
                    6 => std_logic_vector(to_unsigned( 60 , 8)),
                    7 => std_logic_vector(to_unsigned( 9 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=300 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 54 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 83 , 8)),
                    4 => std_logic_vector(to_unsigned( 66 , 8)),
                    5 => std_logic_vector(to_unsigned( 18 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 111 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=301 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 54 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 83 , 8)),
                    4 => std_logic_vector(to_unsigned( 66 , 8)),
                    5 => std_logic_vector(to_unsigned( 18 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 111 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=302 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 112 , 8)),
                    2 => std_logic_vector(to_unsigned( 19 , 8)),
                    3 => std_logic_vector(to_unsigned( 92 , 8)),
                    4 => std_logic_vector(to_unsigned( 116 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 59 , 8)),
                    7 => std_logic_vector(to_unsigned( 79 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=303 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 112 , 8)),
                    4 => std_logic_vector(to_unsigned( 41 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 19 , 8)),
                    7 => std_logic_vector(to_unsigned( 103 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=304 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 112 , 8)),
                    4 => std_logic_vector(to_unsigned( 41 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 19 , 8)),
                    7 => std_logic_vector(to_unsigned( 103 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=305 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 73, 8)),
                    1 => std_logic_vector(to_unsigned( 53 , 8)),
                    2 => std_logic_vector(to_unsigned( 94 , 8)),
                    3 => std_logic_vector(to_unsigned( 116 , 8)),
                    4 => std_logic_vector(to_unsigned( 42 , 8)),
                    5 => std_logic_vector(to_unsigned( 78 , 8)),
                    6 => std_logic_vector(to_unsigned( 17 , 8)),
                    7 => std_logic_vector(to_unsigned( 64 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=306 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 15 , 8)),
                    3 => std_logic_vector(to_unsigned( 106 , 8)),
                    4 => std_logic_vector(to_unsigned( 10 , 8)),
                    5 => std_logic_vector(to_unsigned( 6 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 30 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=307 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 15 , 8)),
                    3 => std_logic_vector(to_unsigned( 106 , 8)),
                    4 => std_logic_vector(to_unsigned( 10 , 8)),
                    5 => std_logic_vector(to_unsigned( 6 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 30 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=308 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),
                    1 => std_logic_vector(to_unsigned( 29 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 19 , 8)),
                    4 => std_logic_vector(to_unsigned( 57 , 8)),
                    5 => std_logic_vector(to_unsigned( 11 , 8)),
                    6 => std_logic_vector(to_unsigned( 61 , 8)),
                    7 => std_logic_vector(to_unsigned( 66 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=309 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 77, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 33 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 21 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=310 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 77, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 33 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 21 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=311 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),
                    1 => std_logic_vector(to_unsigned( 7 , 8)),
                    2 => std_logic_vector(to_unsigned( 73 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 22 , 8)),
                    5 => std_logic_vector(to_unsigned( 124 , 8)),
                    6 => std_logic_vector(to_unsigned( 57 , 8)),
                    7 => std_logic_vector(to_unsigned( 18 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=312 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 40 , 8)),
                    4 => std_logic_vector(to_unsigned( 22 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 83 , 8)),
                    7 => std_logic_vector(to_unsigned( 94 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=313 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 40 , 8)),
                    4 => std_logic_vector(to_unsigned( 22 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 83 , 8)),
                    7 => std_logic_vector(to_unsigned( 94 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=314 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 28 , 8)),
                    3 => std_logic_vector(to_unsigned( 68 , 8)),
                    4 => std_logic_vector(to_unsigned( 49 , 8)),
                    5 => std_logic_vector(to_unsigned( 0 , 8)),
                    6 => std_logic_vector(to_unsigned( 19 , 8)),
                    7 => std_logic_vector(to_unsigned( 96 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=315 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 61 , 8)),
                    2 => std_logic_vector(to_unsigned( 92 , 8)),
                    3 => std_logic_vector(to_unsigned( 23 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 54 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=316 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 61 , 8)),
                    2 => std_logic_vector(to_unsigned( 92 , 8)),
                    3 => std_logic_vector(to_unsigned( 23 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 54 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=317 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 35 , 8)),
                    4 => std_logic_vector(to_unsigned( 98 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 5 , 8)),
                    7 => std_logic_vector(to_unsigned( 48 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=318 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),
                    1 => std_logic_vector(to_unsigned( 96 , 8)),
                    2 => std_logic_vector(to_unsigned( 32 , 8)),
                    3 => std_logic_vector(to_unsigned( 92 , 8)),
                    4 => std_logic_vector(to_unsigned( 67 , 8)),
                    5 => std_logic_vector(to_unsigned( 122 , 8)),
                    6 => std_logic_vector(to_unsigned( 24 , 8)),
                    7 => std_logic_vector(to_unsigned( 82 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=319 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),
                    1 => std_logic_vector(to_unsigned( 96 , 8)),
                    2 => std_logic_vector(to_unsigned( 32 , 8)),
                    3 => std_logic_vector(to_unsigned( 92 , 8)),
                    4 => std_logic_vector(to_unsigned( 67 , 8)),
                    5 => std_logic_vector(to_unsigned( 122 , 8)),
                    6 => std_logic_vector(to_unsigned( 24 , 8)),
                    7 => std_logic_vector(to_unsigned( 82 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=320 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 41, 8)),
                    1 => std_logic_vector(to_unsigned( 101 , 8)),
                    2 => std_logic_vector(to_unsigned( 90 , 8)),
                    3 => std_logic_vector(to_unsigned( 81 , 8)),
                    4 => std_logic_vector(to_unsigned( 2 , 8)),
                    5 => std_logic_vector(to_unsigned( 119 , 8)),
                    6 => std_logic_vector(to_unsigned( 35 , 8)),
                    7 => std_logic_vector(to_unsigned( 94 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=321 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 13 , 8)),
                    4 => std_logic_vector(to_unsigned( 99 , 8)),
                    5 => std_logic_vector(to_unsigned( 8 , 8)),
                    6 => std_logic_vector(to_unsigned( 88 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=322 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 13 , 8)),
                    4 => std_logic_vector(to_unsigned( 99 , 8)),
                    5 => std_logic_vector(to_unsigned( 8 , 8)),
                    6 => std_logic_vector(to_unsigned( 88 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=323 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 82, 8)),
                    1 => std_logic_vector(to_unsigned( 62 , 8)),
                    2 => std_logic_vector(to_unsigned( 86 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 2 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 98 , 8)),
                    7 => std_logic_vector(to_unsigned( 116 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=324 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 49 , 8)),
                    3 => std_logic_vector(to_unsigned( 45 , 8)),
                    4 => std_logic_vector(to_unsigned( 3 , 8)),
                    5 => std_logic_vector(to_unsigned( 24 , 8)),
                    6 => std_logic_vector(to_unsigned( 38 , 8)),
                    7 => std_logic_vector(to_unsigned( 53 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=325 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 49 , 8)),
                    3 => std_logic_vector(to_unsigned( 45 , 8)),
                    4 => std_logic_vector(to_unsigned( 3 , 8)),
                    5 => std_logic_vector(to_unsigned( 24 , 8)),
                    6 => std_logic_vector(to_unsigned( 38 , 8)),
                    7 => std_logic_vector(to_unsigned( 53 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=326 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 27 , 8)),
                    5 => std_logic_vector(to_unsigned( 84 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 33 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=327 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 38 , 8)),
                    2 => std_logic_vector(to_unsigned( 1 , 8)),
                    3 => std_logic_vector(to_unsigned( 105 , 8)),
                    4 => std_logic_vector(to_unsigned( 93 , 8)),
                    5 => std_logic_vector(to_unsigned( 121 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 64 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=328 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 38 , 8)),
                    2 => std_logic_vector(to_unsigned( 1 , 8)),
                    3 => std_logic_vector(to_unsigned( 105 , 8)),
                    4 => std_logic_vector(to_unsigned( 93 , 8)),
                    5 => std_logic_vector(to_unsigned( 121 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 64 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=329 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),
                    1 => std_logic_vector(to_unsigned( 59 , 8)),
                    2 => std_logic_vector(to_unsigned( 29 , 8)),
                    3 => std_logic_vector(to_unsigned( 98 , 8)),
                    4 => std_logic_vector(to_unsigned( 18 , 8)),
                    5 => std_logic_vector(to_unsigned( 111 , 8)),
                    6 => std_logic_vector(to_unsigned( 14 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=330 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 98 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 57 , 8)),
                    4 => std_logic_vector(to_unsigned( 39 , 8)),
                    5 => std_logic_vector(to_unsigned( 13 , 8)),
                    6 => std_logic_vector(to_unsigned( 65 , 8)),
                    7 => std_logic_vector(to_unsigned( 70 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=331 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 98 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 57 , 8)),
                    4 => std_logic_vector(to_unsigned( 39 , 8)),
                    5 => std_logic_vector(to_unsigned( 13 , 8)),
                    6 => std_logic_vector(to_unsigned( 65 , 8)),
                    7 => std_logic_vector(to_unsigned( 70 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=332 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 42, 8)),
                    1 => std_logic_vector(to_unsigned( 17 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 13 , 8)),
                    4 => std_logic_vector(to_unsigned( 22 , 8)),
                    5 => std_logic_vector(to_unsigned( 29 , 8)),
                    6 => std_logic_vector(to_unsigned( 82 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=333 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),
                    1 => std_logic_vector(to_unsigned( 3 , 8)),
                    2 => std_logic_vector(to_unsigned( 20 , 8)),
                    3 => std_logic_vector(to_unsigned( 15 , 8)),
                    4 => std_logic_vector(to_unsigned( 73 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 90 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=334 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),
                    1 => std_logic_vector(to_unsigned( 3 , 8)),
                    2 => std_logic_vector(to_unsigned( 20 , 8)),
                    3 => std_logic_vector(to_unsigned( 15 , 8)),
                    4 => std_logic_vector(to_unsigned( 73 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 90 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=335 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 90, 8)),
                    1 => std_logic_vector(to_unsigned( 77 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 59 , 8)),
                    4 => std_logic_vector(to_unsigned( 9 , 8)),
                    5 => std_logic_vector(to_unsigned( 95 , 8)),
                    6 => std_logic_vector(to_unsigned( 25 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=336 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 57 , 8)),
                    3 => std_logic_vector(to_unsigned( 107 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 15 , 8)),
                    6 => std_logic_vector(to_unsigned( 83 , 8)),
                    7 => std_logic_vector(to_unsigned( 61 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=337 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 57 , 8)),
                    3 => std_logic_vector(to_unsigned( 107 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 15 , 8)),
                    6 => std_logic_vector(to_unsigned( 83 , 8)),
                    7 => std_logic_vector(to_unsigned( 61 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=338 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),
                    1 => std_logic_vector(to_unsigned( 82 , 8)),
                    2 => std_logic_vector(to_unsigned( 31 , 8)),
                    3 => std_logic_vector(to_unsigned( 117 , 8)),
                    4 => std_logic_vector(to_unsigned( 12 , 8)),
                    5 => std_logic_vector(to_unsigned( 2 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=339 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),
                    1 => std_logic_vector(to_unsigned( 57 , 8)),
                    2 => std_logic_vector(to_unsigned( 115 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 75 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 38 , 8)),
                    7 => std_logic_vector(to_unsigned( 12 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=340 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),
                    1 => std_logic_vector(to_unsigned( 57 , 8)),
                    2 => std_logic_vector(to_unsigned( 115 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 75 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 38 , 8)),
                    7 => std_logic_vector(to_unsigned( 12 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=341 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 94 , 8)),
                    2 => std_logic_vector(to_unsigned( 45 , 8)),
                    3 => std_logic_vector(to_unsigned( 8 , 8)),
                    4 => std_logic_vector(to_unsigned( 75 , 8)),
                    5 => std_logic_vector(to_unsigned( 120 , 8)),
                    6 => std_logic_vector(to_unsigned( 1 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=342 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 89 , 8)),
                    2 => std_logic_vector(to_unsigned( 104 , 8)),
                    3 => std_logic_vector(to_unsigned( 56 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 70 , 8)),
                    6 => std_logic_vector(to_unsigned( 79 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=343 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 89 , 8)),
                    2 => std_logic_vector(to_unsigned( 104 , 8)),
                    3 => std_logic_vector(to_unsigned( 56 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 70 , 8)),
                    6 => std_logic_vector(to_unsigned( 79 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=344 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 29 , 8)),
                    2 => std_logic_vector(to_unsigned( 103 , 8)),
                    3 => std_logic_vector(to_unsigned( 5 , 8)),
                    4 => std_logic_vector(to_unsigned( 41 , 8)),
                    5 => std_logic_vector(to_unsigned( 93 , 8)),
                    6 => std_logic_vector(to_unsigned( 35 , 8)),
                    7 => std_logic_vector(to_unsigned( 117 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=345 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 23 , 8)),
                    3 => std_logic_vector(to_unsigned( 71 , 8)),
                    4 => std_logic_vector(to_unsigned( 77 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 104 , 8)),
                    7 => std_logic_vector(to_unsigned( 29 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=346 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 23 , 8)),
                    3 => std_logic_vector(to_unsigned( 71 , 8)),
                    4 => std_logic_vector(to_unsigned( 77 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 104 , 8)),
                    7 => std_logic_vector(to_unsigned( 29 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=347 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 48 , 8)),
                    2 => std_logic_vector(to_unsigned( 81 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 121 , 8)),
                    5 => std_logic_vector(to_unsigned( 77 , 8)),
                    6 => std_logic_vector(to_unsigned( 24 , 8)),
                    7 => std_logic_vector(to_unsigned( 33 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=348 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 53 , 8)),
                    3 => std_logic_vector(to_unsigned( 16 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 118 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=349 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 53 , 8)),
                    3 => std_logic_vector(to_unsigned( 16 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 118 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=350 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 2, 8)),
                    1 => std_logic_vector(to_unsigned( 62 , 8)),
                    2 => std_logic_vector(to_unsigned( 85 , 8)),
                    3 => std_logic_vector(to_unsigned( 116 , 8)),
                    4 => std_logic_vector(to_unsigned( 94 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 48 , 8)),
                    7 => std_logic_vector(to_unsigned( 74 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=351 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 99 , 8)),
                    2 => std_logic_vector(to_unsigned( 122 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 94 , 8)),
                    6 => std_logic_vector(to_unsigned( 78 , 8)),
                    7 => std_logic_vector(to_unsigned( 27 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=352 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 99 , 8)),
                    2 => std_logic_vector(to_unsigned( 122 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 94 , 8)),
                    6 => std_logic_vector(to_unsigned( 78 , 8)),
                    7 => std_logic_vector(to_unsigned( 27 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=353 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 4, 8)),
                    1 => std_logic_vector(to_unsigned( 71 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 43 , 8)),
                    4 => std_logic_vector(to_unsigned( 83 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 15 , 8)),
                    7 => std_logic_vector(to_unsigned( 19 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=354 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 45 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 82 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 123 , 8)),
                    6 => std_logic_vector(to_unsigned( 105 , 8)),
                    7 => std_logic_vector(to_unsigned( 60 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=355 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 45 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 82 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 123 , 8)),
                    6 => std_logic_vector(to_unsigned( 105 , 8)),
                    7 => std_logic_vector(to_unsigned( 60 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=356 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),
                    1 => std_logic_vector(to_unsigned( 15 , 8)),
                    2 => std_logic_vector(to_unsigned( 9 , 8)),
                    3 => std_logic_vector(to_unsigned( 21 , 8)),
                    4 => std_logic_vector(to_unsigned( 30 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 38 , 8)),
                    7 => std_logic_vector(to_unsigned( 112 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=357 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 59 , 8)),
                    3 => std_logic_vector(to_unsigned( 19 , 8)),
                    4 => std_logic_vector(to_unsigned( 26 , 8)),
                    5 => std_logic_vector(to_unsigned( 10 , 8)),
                    6 => std_logic_vector(to_unsigned( 81 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=358 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 59 , 8)),
                    3 => std_logic_vector(to_unsigned( 19 , 8)),
                    4 => std_logic_vector(to_unsigned( 26 , 8)),
                    5 => std_logic_vector(to_unsigned( 10 , 8)),
                    6 => std_logic_vector(to_unsigned( 81 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=359 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 74 , 8)),
                    3 => std_logic_vector(to_unsigned( 57 , 8)),
                    4 => std_logic_vector(to_unsigned( 67 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 14 , 8)),
                    7 => std_logic_vector(to_unsigned( 5 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=360 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),
                    1 => std_logic_vector(to_unsigned( 90 , 8)),
                    2 => std_logic_vector(to_unsigned( 73 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 27 , 8)),
                    5 => std_logic_vector(to_unsigned( 1 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=361 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),
                    1 => std_logic_vector(to_unsigned( 90 , 8)),
                    2 => std_logic_vector(to_unsigned( 73 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 27 , 8)),
                    5 => std_logic_vector(to_unsigned( 1 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=362 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 85 , 8)),
                    3 => std_logic_vector(to_unsigned( 58 , 8)),
                    4 => std_logic_vector(to_unsigned( 22 , 8)),
                    5 => std_logic_vector(to_unsigned( 30 , 8)),
                    6 => std_logic_vector(to_unsigned( 54 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=363 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 50 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 57 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=364 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 50 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 57 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=365 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),
                    1 => std_logic_vector(to_unsigned( 79 , 8)),
                    2 => std_logic_vector(to_unsigned( 58 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 88 , 8)),
                    5 => std_logic_vector(to_unsigned( 6 , 8)),
                    6 => std_logic_vector(to_unsigned( 112 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=366 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 20 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=367 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 20 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=368 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),
                    1 => std_logic_vector(to_unsigned( 92 , 8)),
                    2 => std_logic_vector(to_unsigned( 73 , 8)),
                    3 => std_logic_vector(to_unsigned( 63 , 8)),
                    4 => std_logic_vector(to_unsigned( 118 , 8)),
                    5 => std_logic_vector(to_unsigned( 99 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 57 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=369 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),
                    1 => std_logic_vector(to_unsigned( 65 , 8)),
                    2 => std_logic_vector(to_unsigned( 106 , 8)),
                    3 => std_logic_vector(to_unsigned( 101 , 8)),
                    4 => std_logic_vector(to_unsigned( 121 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 14 , 8)),
                    7 => std_logic_vector(to_unsigned( 42 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=370 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),
                    1 => std_logic_vector(to_unsigned( 65 , 8)),
                    2 => std_logic_vector(to_unsigned( 106 , 8)),
                    3 => std_logic_vector(to_unsigned( 101 , 8)),
                    4 => std_logic_vector(to_unsigned( 121 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 14 , 8)),
                    7 => std_logic_vector(to_unsigned( 42 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=371 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 1 , 8)),
                    3 => std_logic_vector(to_unsigned( 119 , 8)),
                    4 => std_logic_vector(to_unsigned( 38 , 8)),
                    5 => std_logic_vector(to_unsigned( 8 , 8)),
                    6 => std_logic_vector(to_unsigned( 111 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=372 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 114, 8)),
                    1 => std_logic_vector(to_unsigned( 62 , 8)),
                    2 => std_logic_vector(to_unsigned( 99 , 8)),
                    3 => std_logic_vector(to_unsigned( 92 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 68 , 8)),
                    6 => std_logic_vector(to_unsigned( 76 , 8)),
                    7 => std_logic_vector(to_unsigned( 33 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=373 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 114, 8)),
                    1 => std_logic_vector(to_unsigned( 62 , 8)),
                    2 => std_logic_vector(to_unsigned( 99 , 8)),
                    3 => std_logic_vector(to_unsigned( 92 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 68 , 8)),
                    6 => std_logic_vector(to_unsigned( 76 , 8)),
                    7 => std_logic_vector(to_unsigned( 33 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=374 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 96 , 8)),
                    2 => std_logic_vector(to_unsigned( 106 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 43 , 8)),
                    5 => std_logic_vector(to_unsigned( 0 , 8)),
                    6 => std_logic_vector(to_unsigned( 92 , 8)),
                    7 => std_logic_vector(to_unsigned( 16 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=375 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 41 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 28 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=376 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 41 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 28 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=377 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),
                    1 => std_logic_vector(to_unsigned( 93 , 8)),
                    2 => std_logic_vector(to_unsigned( 101 , 8)),
                    3 => std_logic_vector(to_unsigned( 13 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 35 , 8)),
                    7 => std_logic_vector(to_unsigned( 120 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=378 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 14 , 8)),
                    3 => std_logic_vector(to_unsigned( 102 , 8)),
                    4 => std_logic_vector(to_unsigned( 59 , 8)),
                    5 => std_logic_vector(to_unsigned( 55 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 25 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=379 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 14 , 8)),
                    3 => std_logic_vector(to_unsigned( 102 , 8)),
                    4 => std_logic_vector(to_unsigned( 59 , 8)),
                    5 => std_logic_vector(to_unsigned( 55 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 25 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=380 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 113, 8)),
                    1 => std_logic_vector(to_unsigned( 84 , 8)),
                    2 => std_logic_vector(to_unsigned( 43 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 25 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 66 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=381 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 53 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 58 , 8)),
                    4 => std_logic_vector(to_unsigned( 67 , 8)),
                    5 => std_logic_vector(to_unsigned( 101 , 8)),
                    6 => std_logic_vector(to_unsigned( 10 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=382 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 53 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 58 , 8)),
                    4 => std_logic_vector(to_unsigned( 67 , 8)),
                    5 => std_logic_vector(to_unsigned( 101 , 8)),
                    6 => std_logic_vector(to_unsigned( 10 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=383 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),
                    1 => std_logic_vector(to_unsigned( 5 , 8)),
                    2 => std_logic_vector(to_unsigned( 58 , 8)),
                    3 => std_logic_vector(to_unsigned( 67 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 121 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=384 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 38, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 115 , 8)),
                    3 => std_logic_vector(to_unsigned( 62 , 8)),
                    4 => std_logic_vector(to_unsigned( 3 , 8)),
                    5 => std_logic_vector(to_unsigned( 24 , 8)),
                    6 => std_logic_vector(to_unsigned( 19 , 8)),
                    7 => std_logic_vector(to_unsigned( 68 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=385 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 38, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 115 , 8)),
                    3 => std_logic_vector(to_unsigned( 62 , 8)),
                    4 => std_logic_vector(to_unsigned( 3 , 8)),
                    5 => std_logic_vector(to_unsigned( 24 , 8)),
                    6 => std_logic_vector(to_unsigned( 19 , 8)),
                    7 => std_logic_vector(to_unsigned( 68 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=386 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 46, 8)),
                    1 => std_logic_vector(to_unsigned( 20 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 10 , 8)),
                    4 => std_logic_vector(to_unsigned( 79 , 8)),
                    5 => std_logic_vector(to_unsigned( 83 , 8)),
                    6 => std_logic_vector(to_unsigned( 42 , 8)),
                    7 => std_logic_vector(to_unsigned( 25 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=387 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 20 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 112 , 8)),
                    7 => std_logic_vector(to_unsigned( 7 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=388 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 20 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 112 , 8)),
                    7 => std_logic_vector(to_unsigned( 7 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=389 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 52 , 8)),
                    2 => std_logic_vector(to_unsigned( 96 , 8)),
                    3 => std_logic_vector(to_unsigned( 79 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 115 , 8)),
                    6 => std_logic_vector(to_unsigned( 72 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=390 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),
                    1 => std_logic_vector(to_unsigned( 85 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 97 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 109 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=391 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),
                    1 => std_logic_vector(to_unsigned( 85 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 97 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 109 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=392 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 97, 8)),
                    1 => std_logic_vector(to_unsigned( 37 , 8)),
                    2 => std_logic_vector(to_unsigned( 18 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 47 , 8)),
                    5 => std_logic_vector(to_unsigned( 75 , 8)),
                    6 => std_logic_vector(to_unsigned( 14 , 8)),
                    7 => std_logic_vector(to_unsigned( 103 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=393 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 114, 8)),
                    1 => std_logic_vector(to_unsigned( 79 , 8)),
                    2 => std_logic_vector(to_unsigned( 12 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 85 , 8)),
                    5 => std_logic_vector(to_unsigned( 2 , 8)),
                    6 => std_logic_vector(to_unsigned( 49 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=394 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 114, 8)),
                    1 => std_logic_vector(to_unsigned( 79 , 8)),
                    2 => std_logic_vector(to_unsigned( 12 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 85 , 8)),
                    5 => std_logic_vector(to_unsigned( 2 , 8)),
                    6 => std_logic_vector(to_unsigned( 49 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=395 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 60 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 84 , 8)),
                    5 => std_logic_vector(to_unsigned( 5 , 8)),
                    6 => std_logic_vector(to_unsigned( 12 , 8)),
                    7 => std_logic_vector(to_unsigned( 42 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=396 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),
                    1 => std_logic_vector(to_unsigned( 40 , 8)),
                    2 => std_logic_vector(to_unsigned( 65 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 54 , 8)),
                    6 => std_logic_vector(to_unsigned( 69 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=397 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),
                    1 => std_logic_vector(to_unsigned( 40 , 8)),
                    2 => std_logic_vector(to_unsigned( 65 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 54 , 8)),
                    6 => std_logic_vector(to_unsigned( 69 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=398 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),
                    1 => std_logic_vector(to_unsigned( 12 , 8)),
                    2 => std_logic_vector(to_unsigned( 6 , 8)),
                    3 => std_logic_vector(to_unsigned( 119 , 8)),
                    4 => std_logic_vector(to_unsigned( 84 , 8)),
                    5 => std_logic_vector(to_unsigned( 77 , 8)),
                    6 => std_logic_vector(to_unsigned( 44 , 8)),
                    7 => std_logic_vector(to_unsigned( 19 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=399 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 82 , 8)),
                    2 => std_logic_vector(to_unsigned( 46 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 54 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 111 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=400 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 82 , 8)),
                    2 => std_logic_vector(to_unsigned( 46 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 54 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 111 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=401 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 99, 8)),
                    1 => std_logic_vector(to_unsigned( 42 , 8)),
                    2 => std_logic_vector(to_unsigned( 54 , 8)),
                    3 => std_logic_vector(to_unsigned( 92 , 8)),
                    4 => std_logic_vector(to_unsigned( 82 , 8)),
                    5 => std_logic_vector(to_unsigned( 18 , 8)),
                    6 => std_logic_vector(to_unsigned( 29 , 8)),
                    7 => std_logic_vector(to_unsigned( 3 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=402 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 32 , 8)),
                    3 => std_logic_vector(to_unsigned( 109 , 8)),
                    4 => std_logic_vector(to_unsigned( 27 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 60 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=403 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 32 , 8)),
                    3 => std_logic_vector(to_unsigned( 109 , 8)),
                    4 => std_logic_vector(to_unsigned( 27 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 60 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=404 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 100 , 8)),
                    2 => std_logic_vector(to_unsigned( 96 , 8)),
                    3 => std_logic_vector(to_unsigned( 42 , 8)),
                    4 => std_logic_vector(to_unsigned( 82 , 8)),
                    5 => std_logic_vector(to_unsigned( 62 , 8)),
                    6 => std_logic_vector(to_unsigned( 31 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=405 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 2 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 114 , 8)),
                    5 => std_logic_vector(to_unsigned( 55 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=406 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 2 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 114 , 8)),
                    5 => std_logic_vector(to_unsigned( 55 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=407 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),
                    1 => std_logic_vector(to_unsigned( 15 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 123 , 8)),
                    4 => std_logic_vector(to_unsigned( 96 , 8)),
                    5 => std_logic_vector(to_unsigned( 47 , 8)),
                    6 => std_logic_vector(to_unsigned( 82 , 8)),
                    7 => std_logic_vector(to_unsigned( 101 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=408 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 88, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 33 , 8)),
                    6 => std_logic_vector(to_unsigned( 42 , 8)),
                    7 => std_logic_vector(to_unsigned( 15 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=409 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 88, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 33 , 8)),
                    6 => std_logic_vector(to_unsigned( 42 , 8)),
                    7 => std_logic_vector(to_unsigned( 15 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=410 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 44 , 8)),
                    2 => std_logic_vector(to_unsigned( 65 , 8)),
                    3 => std_logic_vector(to_unsigned( 120 , 8)),
                    4 => std_logic_vector(to_unsigned( 33 , 8)),
                    5 => std_logic_vector(to_unsigned( 105 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 14 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=411 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),
                    1 => std_logic_vector(to_unsigned( 53 , 8)),
                    2 => std_logic_vector(to_unsigned( 87 , 8)),
                    3 => std_logic_vector(to_unsigned( 70 , 8)),
                    4 => std_logic_vector(to_unsigned( 124 , 8)),
                    5 => std_logic_vector(to_unsigned( 39 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 110 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=412 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),
                    1 => std_logic_vector(to_unsigned( 53 , 8)),
                    2 => std_logic_vector(to_unsigned( 87 , 8)),
                    3 => std_logic_vector(to_unsigned( 70 , 8)),
                    4 => std_logic_vector(to_unsigned( 124 , 8)),
                    5 => std_logic_vector(to_unsigned( 39 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 110 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=413 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),
                    1 => std_logic_vector(to_unsigned( 53 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 119 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 94 , 8)),
                    6 => std_logic_vector(to_unsigned( 35 , 8)),
                    7 => std_logic_vector(to_unsigned( 74 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=414 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),
                    1 => std_logic_vector(to_unsigned( 80 , 8)),
                    2 => std_logic_vector(to_unsigned( 89 , 8)),
                    3 => std_logic_vector(to_unsigned( 41 , 8)),
                    4 => std_logic_vector(to_unsigned( 105 , 8)),
                    5 => std_logic_vector(to_unsigned( 17 , 8)),
                    6 => std_logic_vector(to_unsigned( 36 , 8)),
                    7 => std_logic_vector(to_unsigned( 9 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=415 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),
                    1 => std_logic_vector(to_unsigned( 80 , 8)),
                    2 => std_logic_vector(to_unsigned( 89 , 8)),
                    3 => std_logic_vector(to_unsigned( 41 , 8)),
                    4 => std_logic_vector(to_unsigned( 105 , 8)),
                    5 => std_logic_vector(to_unsigned( 17 , 8)),
                    6 => std_logic_vector(to_unsigned( 36 , 8)),
                    7 => std_logic_vector(to_unsigned( 9 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=416 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),
                    1 => std_logic_vector(to_unsigned( 29 , 8)),
                    2 => std_logic_vector(to_unsigned( 71 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 114 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 108 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=417 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),
                    1 => std_logic_vector(to_unsigned( 86 , 8)),
                    2 => std_logic_vector(to_unsigned( 80 , 8)),
                    3 => std_logic_vector(to_unsigned( 11 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 124 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=418 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),
                    1 => std_logic_vector(to_unsigned( 86 , 8)),
                    2 => std_logic_vector(to_unsigned( 80 , 8)),
                    3 => std_logic_vector(to_unsigned( 11 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 124 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=419 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 73, 8)),
                    1 => std_logic_vector(to_unsigned( 5 , 8)),
                    2 => std_logic_vector(to_unsigned( 42 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 92 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 30 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=420 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 106 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 46 , 8)),
                    6 => std_logic_vector(to_unsigned( 29 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=421 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 106 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 46 , 8)),
                    6 => std_logic_vector(to_unsigned( 29 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=422 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 105, 8)),
                    1 => std_logic_vector(to_unsigned( 14 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 95 , 8)),
                    4 => std_logic_vector(to_unsigned( 27 , 8)),
                    5 => std_logic_vector(to_unsigned( 73 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 117 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=423 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 29 , 8)),
                    3 => std_logic_vector(to_unsigned( 68 , 8)),
                    4 => std_logic_vector(to_unsigned( 1 , 8)),
                    5 => std_logic_vector(to_unsigned( 118 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 22 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=424 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 29 , 8)),
                    3 => std_logic_vector(to_unsigned( 68 , 8)),
                    4 => std_logic_vector(to_unsigned( 1 , 8)),
                    5 => std_logic_vector(to_unsigned( 118 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 22 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=425 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 94, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 71 , 8)),
                    3 => std_logic_vector(to_unsigned( 31 , 8)),
                    4 => std_logic_vector(to_unsigned( 63 , 8)),
                    5 => std_logic_vector(to_unsigned( 43 , 8)),
                    6 => std_logic_vector(to_unsigned( 67 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=426 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 94, 8)),
                    1 => std_logic_vector(to_unsigned( 58 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 75 , 8)),
                    4 => std_logic_vector(to_unsigned( 10 , 8)),
                    5 => std_logic_vector(to_unsigned( 68 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 36 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=427 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 94, 8)),
                    1 => std_logic_vector(to_unsigned( 58 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 75 , 8)),
                    4 => std_logic_vector(to_unsigned( 10 , 8)),
                    5 => std_logic_vector(to_unsigned( 68 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 36 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=428 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 99, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 108 , 8)),
                    3 => std_logic_vector(to_unsigned( 121 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 70 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=429 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 20 , 8)),
                    2 => std_logic_vector(to_unsigned( 37 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 122 , 8)),
                    5 => std_logic_vector(to_unsigned( 47 , 8)),
                    6 => std_logic_vector(to_unsigned( 115 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=430 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 20 , 8)),
                    2 => std_logic_vector(to_unsigned( 37 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 122 , 8)),
                    5 => std_logic_vector(to_unsigned( 47 , 8)),
                    6 => std_logic_vector(to_unsigned( 115 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=431 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 109, 8)),
                    1 => std_logic_vector(to_unsigned( 44 , 8)),
                    2 => std_logic_vector(to_unsigned( 27 , 8)),
                    3 => std_logic_vector(to_unsigned( 19 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 39 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=432 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 54, 8)),
                    1 => std_logic_vector(to_unsigned( 86 , 8)),
                    2 => std_logic_vector(to_unsigned( 42 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 32 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 97 , 8)),
                    7 => std_logic_vector(to_unsigned( 10 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=433 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 54, 8)),
                    1 => std_logic_vector(to_unsigned( 86 , 8)),
                    2 => std_logic_vector(to_unsigned( 42 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 32 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 97 , 8)),
                    7 => std_logic_vector(to_unsigned( 10 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=434 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 51, 8)),
                    1 => std_logic_vector(to_unsigned( 40 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 114 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 32 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=435 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 106, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 38 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 18 , 8)),
                    5 => std_logic_vector(to_unsigned( 73 , 8)),
                    6 => std_logic_vector(to_unsigned( 68 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=436 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 106, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 38 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 18 , 8)),
                    5 => std_logic_vector(to_unsigned( 73 , 8)),
                    6 => std_logic_vector(to_unsigned( 68 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=437 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 62, 8)),
                    1 => std_logic_vector(to_unsigned( 27 , 8)),
                    2 => std_logic_vector(to_unsigned( 93 , 8)),
                    3 => std_logic_vector(to_unsigned( 110 , 8)),
                    4 => std_logic_vector(to_unsigned( 17 , 8)),
                    5 => std_logic_vector(to_unsigned( 41 , 8)),
                    6 => std_logic_vector(to_unsigned( 82 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=438 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),
                    1 => std_logic_vector(to_unsigned( 18 , 8)),
                    2 => std_logic_vector(to_unsigned( 111 , 8)),
                    3 => std_logic_vector(to_unsigned( 117 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 29 , 8)),
                    6 => std_logic_vector(to_unsigned( 85 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=439 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),
                    1 => std_logic_vector(to_unsigned( 18 , 8)),
                    2 => std_logic_vector(to_unsigned( 111 , 8)),
                    3 => std_logic_vector(to_unsigned( 117 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 29 , 8)),
                    6 => std_logic_vector(to_unsigned( 85 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=440 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),
                    1 => std_logic_vector(to_unsigned( 42 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 96 , 8)),
                    5 => std_logic_vector(to_unsigned( 60 , 8)),
                    6 => std_logic_vector(to_unsigned( 89 , 8)),
                    7 => std_logic_vector(to_unsigned( 74 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=441 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 83 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 56 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 25 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=442 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 83 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 56 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 25 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=443 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 104 , 8)),
                    2 => std_logic_vector(to_unsigned( 121 , 8)),
                    3 => std_logic_vector(to_unsigned( 13 , 8)),
                    4 => std_logic_vector(to_unsigned( 9 , 8)),
                    5 => std_logic_vector(to_unsigned( 34 , 8)),
                    6 => std_logic_vector(to_unsigned( 49 , 8)),
                    7 => std_logic_vector(to_unsigned( 82 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=444 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),
                    1 => std_logic_vector(to_unsigned( 124 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 88 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 102 , 8)),
                    7 => std_logic_vector(to_unsigned( 31 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=445 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),
                    1 => std_logic_vector(to_unsigned( 124 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 88 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 102 , 8)),
                    7 => std_logic_vector(to_unsigned( 31 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=446 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 57 , 8)),
                    3 => std_logic_vector(to_unsigned( 19 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 24 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=447 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 72, 8)),
                    1 => std_logic_vector(to_unsigned( 48 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 85 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 102 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 115 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=448 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 72, 8)),
                    1 => std_logic_vector(to_unsigned( 48 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 85 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 102 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 115 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=449 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 75 , 8)),
                    3 => std_logic_vector(to_unsigned( 67 , 8)),
                    4 => std_logic_vector(to_unsigned( 60 , 8)),
                    5 => std_logic_vector(to_unsigned( 119 , 8)),
                    6 => std_logic_vector(to_unsigned( 30 , 8)),
                    7 => std_logic_vector(to_unsigned( 110 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=450 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),
                    1 => std_logic_vector(to_unsigned( 89 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 84 , 8)),
                    5 => std_logic_vector(to_unsigned( 101 , 8)),
                    6 => std_logic_vector(to_unsigned( 124 , 8)),
                    7 => std_logic_vector(to_unsigned( 20 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=451 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),
                    1 => std_logic_vector(to_unsigned( 89 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 84 , 8)),
                    5 => std_logic_vector(to_unsigned( 101 , 8)),
                    6 => std_logic_vector(to_unsigned( 124 , 8)),
                    7 => std_logic_vector(to_unsigned( 20 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=452 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 53, 8)),
                    1 => std_logic_vector(to_unsigned( 37 , 8)),
                    2 => std_logic_vector(to_unsigned( 117 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 13 , 8)),
                    5 => std_logic_vector(to_unsigned( 46 , 8)),
                    6 => std_logic_vector(to_unsigned( 68 , 8)),
                    7 => std_logic_vector(to_unsigned( 103 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=453 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 43 , 8)),
                    5 => std_logic_vector(to_unsigned( 1 , 8)),
                    6 => std_logic_vector(to_unsigned( 33 , 8)),
                    7 => std_logic_vector(to_unsigned( 104 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=454 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 43 , 8)),
                    5 => std_logic_vector(to_unsigned( 1 , 8)),
                    6 => std_logic_vector(to_unsigned( 33 , 8)),
                    7 => std_logic_vector(to_unsigned( 104 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=455 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 94, 8)),
                    1 => std_logic_vector(to_unsigned( 44 , 8)),
                    2 => std_logic_vector(to_unsigned( 59 , 8)),
                    3 => std_logic_vector(to_unsigned( 115 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 2 , 8)),
                    6 => std_logic_vector(to_unsigned( 124 , 8)),
                    7 => std_logic_vector(to_unsigned( 101 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=456 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 62, 8)),
                    1 => std_logic_vector(to_unsigned( 39 , 8)),
                    2 => std_logic_vector(to_unsigned( 113 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 22 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=457 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 62, 8)),
                    1 => std_logic_vector(to_unsigned( 39 , 8)),
                    2 => std_logic_vector(to_unsigned( 113 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 22 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=458 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 63, 8)),
                    1 => std_logic_vector(to_unsigned( 46 , 8)),
                    2 => std_logic_vector(to_unsigned( 30 , 8)),
                    3 => std_logic_vector(to_unsigned( 79 , 8)),
                    4 => std_logic_vector(to_unsigned( 67 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 17 , 8)),
                    7 => std_logic_vector(to_unsigned( 115 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=459 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 4, 8)),
                    1 => std_logic_vector(to_unsigned( 44 , 8)),
                    2 => std_logic_vector(to_unsigned( 98 , 8)),
                    3 => std_logic_vector(to_unsigned( 69 , 8)),
                    4 => std_logic_vector(to_unsigned( 20 , 8)),
                    5 => std_logic_vector(to_unsigned( 93 , 8)),
                    6 => std_logic_vector(to_unsigned( 107 , 8)),
                    7 => std_logic_vector(to_unsigned( 24 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=460 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 4, 8)),
                    1 => std_logic_vector(to_unsigned( 44 , 8)),
                    2 => std_logic_vector(to_unsigned( 98 , 8)),
                    3 => std_logic_vector(to_unsigned( 69 , 8)),
                    4 => std_logic_vector(to_unsigned( 20 , 8)),
                    5 => std_logic_vector(to_unsigned( 93 , 8)),
                    6 => std_logic_vector(to_unsigned( 107 , 8)),
                    7 => std_logic_vector(to_unsigned( 24 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=461 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),
                    1 => std_logic_vector(to_unsigned( 117 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 93 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 73 , 8)),
                    6 => std_logic_vector(to_unsigned( 54 , 8)),
                    7 => std_logic_vector(to_unsigned( 77 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=462 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 71, 8)),
                    1 => std_logic_vector(to_unsigned( 32 , 8)),
                    2 => std_logic_vector(to_unsigned( 47 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 66 , 8)),
                    5 => std_logic_vector(to_unsigned( 110 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 5 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=463 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 71, 8)),
                    1 => std_logic_vector(to_unsigned( 32 , 8)),
                    2 => std_logic_vector(to_unsigned( 47 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 66 , 8)),
                    5 => std_logic_vector(to_unsigned( 110 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 5 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=464 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 9 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 65 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 109 , 8)),
                    7 => std_logic_vector(to_unsigned( 52 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=465 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 105, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 47 , 8)),
                    3 => std_logic_vector(to_unsigned( 14 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 41 , 8)),
                    6 => std_logic_vector(to_unsigned( 10 , 8)),
                    7 => std_logic_vector(to_unsigned( 4 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=466 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 105, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 47 , 8)),
                    3 => std_logic_vector(to_unsigned( 14 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 41 , 8)),
                    6 => std_logic_vector(to_unsigned( 10 , 8)),
                    7 => std_logic_vector(to_unsigned( 4 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=467 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 12 , 8)),
                    2 => std_logic_vector(to_unsigned( 61 , 8)),
                    3 => std_logic_vector(to_unsigned( 86 , 8)),
                    4 => std_logic_vector(to_unsigned( 104 , 8)),
                    5 => std_logic_vector(to_unsigned( 0 , 8)),
                    6 => std_logic_vector(to_unsigned( 114 , 8)),
                    7 => std_logic_vector(to_unsigned( 38 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=468 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),
                    1 => std_logic_vector(to_unsigned( 5 , 8)),
                    2 => std_logic_vector(to_unsigned( 114 , 8)),
                    3 => std_logic_vector(to_unsigned( 70 , 8)),
                    4 => std_logic_vector(to_unsigned( 120 , 8)),
                    5 => std_logic_vector(to_unsigned( 77 , 8)),
                    6 => std_logic_vector(to_unsigned( 30 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=469 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),
                    1 => std_logic_vector(to_unsigned( 5 , 8)),
                    2 => std_logic_vector(to_unsigned( 114 , 8)),
                    3 => std_logic_vector(to_unsigned( 70 , 8)),
                    4 => std_logic_vector(to_unsigned( 120 , 8)),
                    5 => std_logic_vector(to_unsigned( 77 , 8)),
                    6 => std_logic_vector(to_unsigned( 30 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=470 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 89 , 8)),
                    3 => std_logic_vector(to_unsigned( 36 , 8)),
                    4 => std_logic_vector(to_unsigned( 44 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 30 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=471 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),
                    1 => std_logic_vector(to_unsigned( 113 , 8)),
                    2 => std_logic_vector(to_unsigned( 38 , 8)),
                    3 => std_logic_vector(to_unsigned( 75 , 8)),
                    4 => std_logic_vector(to_unsigned( 106 , 8)),
                    5 => std_logic_vector(to_unsigned( 48 , 8)),
                    6 => std_logic_vector(to_unsigned( 32 , 8)),
                    7 => std_logic_vector(to_unsigned( 99 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=472 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),
                    1 => std_logic_vector(to_unsigned( 113 , 8)),
                    2 => std_logic_vector(to_unsigned( 38 , 8)),
                    3 => std_logic_vector(to_unsigned( 75 , 8)),
                    4 => std_logic_vector(to_unsigned( 106 , 8)),
                    5 => std_logic_vector(to_unsigned( 48 , 8)),
                    6 => std_logic_vector(to_unsigned( 32 , 8)),
                    7 => std_logic_vector(to_unsigned( 99 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=473 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 40 , 8)),
                    2 => std_logic_vector(to_unsigned( 50 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 77 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 69 , 8)),
                    7 => std_logic_vector(to_unsigned( 29 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=474 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 3 , 8)),
                    3 => std_logic_vector(to_unsigned( 105 , 8)),
                    4 => std_logic_vector(to_unsigned( 93 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 55 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=475 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 3 , 8)),
                    3 => std_logic_vector(to_unsigned( 105 , 8)),
                    4 => std_logic_vector(to_unsigned( 93 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 55 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=476 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 70 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 111 , 8)),
                    6 => std_logic_vector(to_unsigned( 88 , 8)),
                    7 => std_logic_vector(to_unsigned( 11 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=477 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 120 , 8)),
                    2 => std_logic_vector(to_unsigned( 84 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 97 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 55 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=478 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 120 , 8)),
                    2 => std_logic_vector(to_unsigned( 84 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 97 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 55 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=479 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),
                    1 => std_logic_vector(to_unsigned( 33 , 8)),
                    2 => std_logic_vector(to_unsigned( 78 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 59 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 65 , 8)),
                    7 => std_logic_vector(to_unsigned( 71 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=480 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 71, 8)),
                    1 => std_logic_vector(to_unsigned( 112 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 82 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 22 , 8)),
                    6 => std_logic_vector(to_unsigned( 41 , 8)),
                    7 => std_logic_vector(to_unsigned( 26 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=481 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 71, 8)),
                    1 => std_logic_vector(to_unsigned( 112 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 82 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 22 , 8)),
                    6 => std_logic_vector(to_unsigned( 41 , 8)),
                    7 => std_logic_vector(to_unsigned( 26 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=482 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 114 , 8)),
                    5 => std_logic_vector(to_unsigned( 70 , 8)),
                    6 => std_logic_vector(to_unsigned( 3 , 8)),
                    7 => std_logic_vector(to_unsigned( 77 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=483 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 67, 8)),
                    1 => std_logic_vector(to_unsigned( 111 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 75 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 51 , 8)),
                    6 => std_logic_vector(to_unsigned( 89 , 8)),
                    7 => std_logic_vector(to_unsigned( 57 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=484 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 67, 8)),
                    1 => std_logic_vector(to_unsigned( 111 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 75 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 51 , 8)),
                    6 => std_logic_vector(to_unsigned( 89 , 8)),
                    7 => std_logic_vector(to_unsigned( 57 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=485 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),
                    1 => std_logic_vector(to_unsigned( 45 , 8)),
                    2 => std_logic_vector(to_unsigned( 99 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 80 , 8)),
                    5 => std_logic_vector(to_unsigned( 6 , 8)),
                    6 => std_logic_vector(to_unsigned( 14 , 8)),
                    7 => std_logic_vector(to_unsigned( 70 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=486 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 23 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 102 , 8)),
                    7 => std_logic_vector(to_unsigned( 115 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=487 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 23 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 102 , 8)),
                    7 => std_logic_vector(to_unsigned( 115 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=488 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 70 , 8)),
                    2 => std_logic_vector(to_unsigned( 49 , 8)),
                    3 => std_logic_vector(to_unsigned( 56 , 8)),
                    4 => std_logic_vector(to_unsigned( 31 , 8)),
                    5 => std_logic_vector(to_unsigned( 91 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 19 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=489 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 70 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 33 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=490 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 70 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 33 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=491 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 33 , 8)),
                    2 => std_logic_vector(to_unsigned( 6 , 8)),
                    3 => std_logic_vector(to_unsigned( 2 , 8)),
                    4 => std_logic_vector(to_unsigned( 123 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 113 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=492 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 39, 8)),
                    1 => std_logic_vector(to_unsigned( 14 , 8)),
                    2 => std_logic_vector(to_unsigned( 70 , 8)),
                    3 => std_logic_vector(to_unsigned( 53 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 49 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 64 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=493 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 39, 8)),
                    1 => std_logic_vector(to_unsigned( 14 , 8)),
                    2 => std_logic_vector(to_unsigned( 70 , 8)),
                    3 => std_logic_vector(to_unsigned( 53 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 49 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 64 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=494 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),
                    1 => std_logic_vector(to_unsigned( 105 , 8)),
                    2 => std_logic_vector(to_unsigned( 11 , 8)),
                    3 => std_logic_vector(to_unsigned( 37 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 118 , 8)),
                    6 => std_logic_vector(to_unsigned( 124 , 8)),
                    7 => std_logic_vector(to_unsigned( 22 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=495 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 108 , 8)),
                    3 => std_logic_vector(to_unsigned( 25 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 88 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=496 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 108 , 8)),
                    3 => std_logic_vector(to_unsigned( 25 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 88 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=497 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 2 , 8)),
                    2 => std_logic_vector(to_unsigned( 35 , 8)),
                    3 => std_logic_vector(to_unsigned( 101 , 8)),
                    4 => std_logic_vector(to_unsigned( 14 , 8)),
                    5 => std_logic_vector(to_unsigned( 60 , 8)),
                    6 => std_logic_vector(to_unsigned( 83 , 8)),
                    7 => std_logic_vector(to_unsigned( 19 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=498 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 103 , 8)),
                    2 => std_logic_vector(to_unsigned( 19 , 8)),
                    3 => std_logic_vector(to_unsigned( 118 , 8)),
                    4 => std_logic_vector(to_unsigned( 6 , 8)),
                    5 => std_logic_vector(to_unsigned( 13 , 8)),
                    6 => std_logic_vector(to_unsigned( 124 , 8)),
                    7 => std_logic_vector(to_unsigned( 107 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=499 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 103 , 8)),
                    2 => std_logic_vector(to_unsigned( 19 , 8)),
                    3 => std_logic_vector(to_unsigned( 118 , 8)),
                    4 => std_logic_vector(to_unsigned( 6 , 8)),
                    5 => std_logic_vector(to_unsigned( 13 , 8)),
                    6 => std_logic_vector(to_unsigned( 124 , 8)),
                    7 => std_logic_vector(to_unsigned( 107 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=500 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),
                    1 => std_logic_vector(to_unsigned( 71 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 45 , 8)),
                    4 => std_logic_vector(to_unsigned( 49 , 8)),
                    5 => std_logic_vector(to_unsigned( 82 , 8)),
                    6 => std_logic_vector(to_unsigned( 29 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=501 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),
                    1 => std_logic_vector(to_unsigned( 108 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 34 , 8)),
                    5 => std_logic_vector(to_unsigned( 60 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 52 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=502 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),
                    1 => std_logic_vector(to_unsigned( 108 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 34 , 8)),
                    5 => std_logic_vector(to_unsigned( 60 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 52 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=503 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 65, 8)),
                    1 => std_logic_vector(to_unsigned( 70 , 8)),
                    2 => std_logic_vector(to_unsigned( 86 , 8)),
                    3 => std_logic_vector(to_unsigned( 21 , 8)),
                    4 => std_logic_vector(to_unsigned( 75 , 8)),
                    5 => std_logic_vector(to_unsigned( 91 , 8)),
                    6 => std_logic_vector(to_unsigned( 114 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=504 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 86 , 8)),
                    3 => std_logic_vector(to_unsigned( 50 , 8)),
                    4 => std_logic_vector(to_unsigned( 30 , 8)),
                    5 => std_logic_vector(to_unsigned( 116 , 8)),
                    6 => std_logic_vector(to_unsigned( 15 , 8)),
                    7 => std_logic_vector(to_unsigned( 4 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=505 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 86 , 8)),
                    3 => std_logic_vector(to_unsigned( 50 , 8)),
                    4 => std_logic_vector(to_unsigned( 30 , 8)),
                    5 => std_logic_vector(to_unsigned( 116 , 8)),
                    6 => std_logic_vector(to_unsigned( 15 , 8)),
                    7 => std_logic_vector(to_unsigned( 4 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=506 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 80 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 23 , 8)),
                    6 => std_logic_vector(to_unsigned( 41 , 8)),
                    7 => std_logic_vector(to_unsigned( 120 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=507 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 19 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 48 , 8)),
                    5 => std_logic_vector(to_unsigned( 32 , 8)),
                    6 => std_logic_vector(to_unsigned( 63 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=508 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 19 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 48 , 8)),
                    5 => std_logic_vector(to_unsigned( 32 , 8)),
                    6 => std_logic_vector(to_unsigned( 63 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=509 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 113, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 19 , 8)),
                    3 => std_logic_vector(to_unsigned( 88 , 8)),
                    4 => std_logic_vector(to_unsigned( 38 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 121 , 8)),
                    7 => std_logic_vector(to_unsigned( 29 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=510 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 9, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 91 , 8)),
                    3 => std_logic_vector(to_unsigned( 79 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 99 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=511 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 9, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 91 , 8)),
                    3 => std_logic_vector(to_unsigned( 79 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 99 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=512 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 63, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 45 , 8)),
                    3 => std_logic_vector(to_unsigned( 119 , 8)),
                    4 => std_logic_vector(to_unsigned( 11 , 8)),
                    5 => std_logic_vector(to_unsigned( 90 , 8)),
                    6 => std_logic_vector(to_unsigned( 69 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=513 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 20 , 8)),
                    3 => std_logic_vector(to_unsigned( 107 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=514 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 20 , 8)),
                    3 => std_logic_vector(to_unsigned( 107 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=515 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 113, 8)),
                    1 => std_logic_vector(to_unsigned( 47 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 109 , 8)),
                    6 => std_logic_vector(to_unsigned( 12 , 8)),
                    7 => std_logic_vector(to_unsigned( 54 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=516 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 56 , 8)),
                    4 => std_logic_vector(to_unsigned( 79 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 27 , 8)),
                    7 => std_logic_vector(to_unsigned( 15 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=517 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 56 , 8)),
                    4 => std_logic_vector(to_unsigned( 79 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 27 , 8)),
                    7 => std_logic_vector(to_unsigned( 15 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=518 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 13 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 78 , 8)),
                    5 => std_logic_vector(to_unsigned( 20 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 36 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=519 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 14 , 8)),
                    5 => std_logic_vector(to_unsigned( 10 , 8)),
                    6 => std_logic_vector(to_unsigned( 109 , 8)),
                    7 => std_logic_vector(to_unsigned( 31 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=520 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 14 , 8)),
                    5 => std_logic_vector(to_unsigned( 10 , 8)),
                    6 => std_logic_vector(to_unsigned( 109 , 8)),
                    7 => std_logic_vector(to_unsigned( 31 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=521 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),
                    1 => std_logic_vector(to_unsigned( 82 , 8)),
                    2 => std_logic_vector(to_unsigned( 15 , 8)),
                    3 => std_logic_vector(to_unsigned( 6 , 8)),
                    4 => std_logic_vector(to_unsigned( 54 , 8)),
                    5 => std_logic_vector(to_unsigned( 110 , 8)),
                    6 => std_logic_vector(to_unsigned( 87 , 8)),
                    7 => std_logic_vector(to_unsigned( 48 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=522 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 45 , 8)),
                    2 => std_logic_vector(to_unsigned( 3 , 8)),
                    3 => std_logic_vector(to_unsigned( 18 , 8)),
                    4 => std_logic_vector(to_unsigned( 37 , 8)),
                    5 => std_logic_vector(to_unsigned( 105 , 8)),
                    6 => std_logic_vector(to_unsigned( 65 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=523 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 45 , 8)),
                    2 => std_logic_vector(to_unsigned( 3 , 8)),
                    3 => std_logic_vector(to_unsigned( 18 , 8)),
                    4 => std_logic_vector(to_unsigned( 37 , 8)),
                    5 => std_logic_vector(to_unsigned( 105 , 8)),
                    6 => std_logic_vector(to_unsigned( 65 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=524 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),
                    1 => std_logic_vector(to_unsigned( 7 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 29 , 8)),
                    4 => std_logic_vector(to_unsigned( 17 , 8)),
                    5 => std_logic_vector(to_unsigned( 50 , 8)),
                    6 => std_logic_vector(to_unsigned( 64 , 8)),
                    7 => std_logic_vector(to_unsigned( 55 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=525 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 84, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 97 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 10 , 8)),
                    7 => std_logic_vector(to_unsigned( 52 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=526 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 84, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 97 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 10 , 8)),
                    7 => std_logic_vector(to_unsigned( 52 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=527 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 6 , 8)),
                    3 => std_logic_vector(to_unsigned( 26 , 8)),
                    4 => std_logic_vector(to_unsigned( 98 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 46 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=528 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),
                    1 => std_logic_vector(to_unsigned( 56 , 8)),
                    2 => std_logic_vector(to_unsigned( 14 , 8)),
                    3 => std_logic_vector(to_unsigned( 102 , 8)),
                    4 => std_logic_vector(to_unsigned( 77 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 89 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=529 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),
                    1 => std_logic_vector(to_unsigned( 56 , 8)),
                    2 => std_logic_vector(to_unsigned( 14 , 8)),
                    3 => std_logic_vector(to_unsigned( 102 , 8)),
                    4 => std_logic_vector(to_unsigned( 77 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 89 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=530 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 24 , 8)),
                    3 => std_logic_vector(to_unsigned( 92 , 8)),
                    4 => std_logic_vector(to_unsigned( 6 , 8)),
                    5 => std_logic_vector(to_unsigned( 78 , 8)),
                    6 => std_logic_vector(to_unsigned( 15 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=531 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),
                    1 => std_logic_vector(to_unsigned( 18 , 8)),
                    2 => std_logic_vector(to_unsigned( 59 , 8)),
                    3 => std_logic_vector(to_unsigned( 109 , 8)),
                    4 => std_logic_vector(to_unsigned( 79 , 8)),
                    5 => std_logic_vector(to_unsigned( 94 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 121 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=532 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),
                    1 => std_logic_vector(to_unsigned( 18 , 8)),
                    2 => std_logic_vector(to_unsigned( 59 , 8)),
                    3 => std_logic_vector(to_unsigned( 109 , 8)),
                    4 => std_logic_vector(to_unsigned( 79 , 8)),
                    5 => std_logic_vector(to_unsigned( 94 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 121 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=533 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 84, 8)),
                    1 => std_logic_vector(to_unsigned( 66 , 8)),
                    2 => std_logic_vector(to_unsigned( 74 , 8)),
                    3 => std_logic_vector(to_unsigned( 89 , 8)),
                    4 => std_logic_vector(to_unsigned( 51 , 8)),
                    5 => std_logic_vector(to_unsigned( 27 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 122 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=534 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 96 , 8)),
                    3 => std_logic_vector(to_unsigned( 86 , 8)),
                    4 => std_logic_vector(to_unsigned( 78 , 8)),
                    5 => std_logic_vector(to_unsigned( 10 , 8)),
                    6 => std_logic_vector(to_unsigned( 90 , 8)),
                    7 => std_logic_vector(to_unsigned( 74 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=535 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 96 , 8)),
                    3 => std_logic_vector(to_unsigned( 86 , 8)),
                    4 => std_logic_vector(to_unsigned( 78 , 8)),
                    5 => std_logic_vector(to_unsigned( 10 , 8)),
                    6 => std_logic_vector(to_unsigned( 90 , 8)),
                    7 => std_logic_vector(to_unsigned( 74 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=536 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 42 , 8)),
                    2 => std_logic_vector(to_unsigned( 68 , 8)),
                    3 => std_logic_vector(to_unsigned( 76 , 8)),
                    4 => std_logic_vector(to_unsigned( 37 , 8)),
                    5 => std_logic_vector(to_unsigned( 3 , 8)),
                    6 => std_logic_vector(to_unsigned( 49 , 8)),
                    7 => std_logic_vector(to_unsigned( 113 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=537 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 51, 8)),
                    1 => std_logic_vector(to_unsigned( 124 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 88 , 8)),
                    4 => std_logic_vector(to_unsigned( 39 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 99 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=538 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 51, 8)),
                    1 => std_logic_vector(to_unsigned( 124 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 88 , 8)),
                    4 => std_logic_vector(to_unsigned( 39 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 99 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=539 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 26 , 8)),
                    2 => std_logic_vector(to_unsigned( 103 , 8)),
                    3 => std_logic_vector(to_unsigned( 21 , 8)),
                    4 => std_logic_vector(to_unsigned( 83 , 8)),
                    5 => std_logic_vector(to_unsigned( 87 , 8)),
                    6 => std_logic_vector(to_unsigned( 109 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=540 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 77, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 103 , 8)),
                    4 => std_logic_vector(to_unsigned( 68 , 8)),
                    5 => std_logic_vector(to_unsigned( 12 , 8)),
                    6 => std_logic_vector(to_unsigned( 4 , 8)),
                    7 => std_logic_vector(to_unsigned( 118 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=541 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 77, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 103 , 8)),
                    4 => std_logic_vector(to_unsigned( 68 , 8)),
                    5 => std_logic_vector(to_unsigned( 12 , 8)),
                    6 => std_logic_vector(to_unsigned( 4 , 8)),
                    7 => std_logic_vector(to_unsigned( 118 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=542 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),
                    1 => std_logic_vector(to_unsigned( 124 , 8)),
                    2 => std_logic_vector(to_unsigned( 33 , 8)),
                    3 => std_logic_vector(to_unsigned( 81 , 8)),
                    4 => std_logic_vector(to_unsigned( 13 , 8)),
                    5 => std_logic_vector(to_unsigned( 19 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=543 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),
                    1 => std_logic_vector(to_unsigned( 119 , 8)),
                    2 => std_logic_vector(to_unsigned( 86 , 8)),
                    3 => std_logic_vector(to_unsigned( 18 , 8)),
                    4 => std_logic_vector(to_unsigned( 124 , 8)),
                    5 => std_logic_vector(to_unsigned( 75 , 8)),
                    6 => std_logic_vector(to_unsigned( 46 , 8)),
                    7 => std_logic_vector(to_unsigned( 11 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=544 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),
                    1 => std_logic_vector(to_unsigned( 119 , 8)),
                    2 => std_logic_vector(to_unsigned( 86 , 8)),
                    3 => std_logic_vector(to_unsigned( 18 , 8)),
                    4 => std_logic_vector(to_unsigned( 124 , 8)),
                    5 => std_logic_vector(to_unsigned( 75 , 8)),
                    6 => std_logic_vector(to_unsigned( 46 , 8)),
                    7 => std_logic_vector(to_unsigned( 11 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=545 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),
                    1 => std_logic_vector(to_unsigned( 19 , 8)),
                    2 => std_logic_vector(to_unsigned( 121 , 8)),
                    3 => std_logic_vector(to_unsigned( 43 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 76 , 8)),
                    6 => std_logic_vector(to_unsigned( 54 , 8)),
                    7 => std_logic_vector(to_unsigned( 28 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=546 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 63, 8)),
                    1 => std_logic_vector(to_unsigned( 110 , 8)),
                    2 => std_logic_vector(to_unsigned( 51 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 42 , 8)),
                    5 => std_logic_vector(to_unsigned( 100 , 8)),
                    6 => std_logic_vector(to_unsigned( 22 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=547 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 63, 8)),
                    1 => std_logic_vector(to_unsigned( 110 , 8)),
                    2 => std_logic_vector(to_unsigned( 51 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 42 , 8)),
                    5 => std_logic_vector(to_unsigned( 100 , 8)),
                    6 => std_logic_vector(to_unsigned( 22 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=548 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 54 , 8)),
                    2 => std_logic_vector(to_unsigned( 108 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 29 , 8)),
                    6 => std_logic_vector(to_unsigned( 22 , 8)),
                    7 => std_logic_vector(to_unsigned( 44 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=549 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 84 , 8)),
                    2 => std_logic_vector(to_unsigned( 48 , 8)),
                    3 => std_logic_vector(to_unsigned( 97 , 8)),
                    4 => std_logic_vector(to_unsigned( 43 , 8)),
                    5 => std_logic_vector(to_unsigned( 62 , 8)),
                    6 => std_logic_vector(to_unsigned( 3 , 8)),
                    7 => std_logic_vector(to_unsigned( 74 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=550 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 84 , 8)),
                    2 => std_logic_vector(to_unsigned( 48 , 8)),
                    3 => std_logic_vector(to_unsigned( 97 , 8)),
                    4 => std_logic_vector(to_unsigned( 43 , 8)),
                    5 => std_logic_vector(to_unsigned( 62 , 8)),
                    6 => std_logic_vector(to_unsigned( 3 , 8)),
                    7 => std_logic_vector(to_unsigned( 74 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=551 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),
                    1 => std_logic_vector(to_unsigned( 44 , 8)),
                    2 => std_logic_vector(to_unsigned( 2 , 8)),
                    3 => std_logic_vector(to_unsigned( 122 , 8)),
                    4 => std_logic_vector(to_unsigned( 99 , 8)),
                    5 => std_logic_vector(to_unsigned( 51 , 8)),
                    6 => std_logic_vector(to_unsigned( 81 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=552 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 25, 8)),
                    1 => std_logic_vector(to_unsigned( 56 , 8)),
                    2 => std_logic_vector(to_unsigned( 82 , 8)),
                    3 => std_logic_vector(to_unsigned( 11 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 7 , 8)),
                    6 => std_logic_vector(to_unsigned( 77 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=553 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 25, 8)),
                    1 => std_logic_vector(to_unsigned( 56 , 8)),
                    2 => std_logic_vector(to_unsigned( 82 , 8)),
                    3 => std_logic_vector(to_unsigned( 11 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 7 , 8)),
                    6 => std_logic_vector(to_unsigned( 77 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=554 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 105 , 8)),
                    2 => std_logic_vector(to_unsigned( 12 , 8)),
                    3 => std_logic_vector(to_unsigned( 79 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 64 , 8)),
                    6 => std_logic_vector(to_unsigned( 83 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=555 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 18 , 8)),
                    2 => std_logic_vector(to_unsigned( 56 , 8)),
                    3 => std_logic_vector(to_unsigned( 82 , 8)),
                    4 => std_logic_vector(to_unsigned( 49 , 8)),
                    5 => std_logic_vector(to_unsigned( 71 , 8)),
                    6 => std_logic_vector(to_unsigned( 27 , 8)),
                    7 => std_logic_vector(to_unsigned( 10 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=556 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 18 , 8)),
                    2 => std_logic_vector(to_unsigned( 56 , 8)),
                    3 => std_logic_vector(to_unsigned( 82 , 8)),
                    4 => std_logic_vector(to_unsigned( 49 , 8)),
                    5 => std_logic_vector(to_unsigned( 71 , 8)),
                    6 => std_logic_vector(to_unsigned( 27 , 8)),
                    7 => std_logic_vector(to_unsigned( 10 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=557 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 104 , 8)),
                    2 => std_logic_vector(to_unsigned( 26 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 110 , 8)),
                    5 => std_logic_vector(to_unsigned( 83 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=558 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 17, 8)),
                    1 => std_logic_vector(to_unsigned( 101 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 57 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 91 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 1 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=559 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 17, 8)),
                    1 => std_logic_vector(to_unsigned( 101 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 57 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 91 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 1 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=560 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),
                    1 => std_logic_vector(to_unsigned( 107 , 8)),
                    2 => std_logic_vector(to_unsigned( 56 , 8)),
                    3 => std_logic_vector(to_unsigned( 91 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 75 , 8)),
                    6 => std_logic_vector(to_unsigned( 27 , 8)),
                    7 => std_logic_vector(to_unsigned( 22 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=561 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),
                    1 => std_logic_vector(to_unsigned( 90 , 8)),
                    2 => std_logic_vector(to_unsigned( 11 , 8)),
                    3 => std_logic_vector(to_unsigned( 122 , 8)),
                    4 => std_logic_vector(to_unsigned( 34 , 8)),
                    5 => std_logic_vector(to_unsigned( 29 , 8)),
                    6 => std_logic_vector(to_unsigned( 23 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=562 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),
                    1 => std_logic_vector(to_unsigned( 90 , 8)),
                    2 => std_logic_vector(to_unsigned( 11 , 8)),
                    3 => std_logic_vector(to_unsigned( 122 , 8)),
                    4 => std_logic_vector(to_unsigned( 34 , 8)),
                    5 => std_logic_vector(to_unsigned( 29 , 8)),
                    6 => std_logic_vector(to_unsigned( 23 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=563 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 120 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 97 , 8)),
                    5 => std_logic_vector(to_unsigned( 115 , 8)),
                    6 => std_logic_vector(to_unsigned( 107 , 8)),
                    7 => std_logic_vector(to_unsigned( 18 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=564 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),
                    1 => std_logic_vector(to_unsigned( 98 , 8)),
                    2 => std_logic_vector(to_unsigned( 105 , 8)),
                    3 => std_logic_vector(to_unsigned( 76 , 8)),
                    4 => std_logic_vector(to_unsigned( 87 , 8)),
                    5 => std_logic_vector(to_unsigned( 82 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 113 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=565 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),
                    1 => std_logic_vector(to_unsigned( 98 , 8)),
                    2 => std_logic_vector(to_unsigned( 105 , 8)),
                    3 => std_logic_vector(to_unsigned( 76 , 8)),
                    4 => std_logic_vector(to_unsigned( 87 , 8)),
                    5 => std_logic_vector(to_unsigned( 82 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 113 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=566 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 39 , 8)),
                    2 => std_logic_vector(to_unsigned( 117 , 8)),
                    3 => std_logic_vector(to_unsigned( 27 , 8)),
                    4 => std_logic_vector(to_unsigned( 96 , 8)),
                    5 => std_logic_vector(to_unsigned( 18 , 8)),
                    6 => std_logic_vector(to_unsigned( 8 , 8)),
                    7 => std_logic_vector(to_unsigned( 113 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=567 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),
                    1 => std_logic_vector(to_unsigned( 16 , 8)),
                    2 => std_logic_vector(to_unsigned( 37 , 8)),
                    3 => std_logic_vector(to_unsigned( 60 , 8)),
                    4 => std_logic_vector(to_unsigned( 49 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 20 , 8)),
                    7 => std_logic_vector(to_unsigned( 27 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=568 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),
                    1 => std_logic_vector(to_unsigned( 16 , 8)),
                    2 => std_logic_vector(to_unsigned( 37 , 8)),
                    3 => std_logic_vector(to_unsigned( 60 , 8)),
                    4 => std_logic_vector(to_unsigned( 49 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 20 , 8)),
                    7 => std_logic_vector(to_unsigned( 27 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=569 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),
                    1 => std_logic_vector(to_unsigned( 48 , 8)),
                    2 => std_logic_vector(to_unsigned( 98 , 8)),
                    3 => std_logic_vector(to_unsigned( 67 , 8)),
                    4 => std_logic_vector(to_unsigned( 105 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 42 , 8)),
                    7 => std_logic_vector(to_unsigned( 90 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=570 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 80, 8)),
                    1 => std_logic_vector(to_unsigned( 37 , 8)),
                    2 => std_logic_vector(to_unsigned( 100 , 8)),
                    3 => std_logic_vector(to_unsigned( 2 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 93 , 8)),
                    6 => std_logic_vector(to_unsigned( 52 , 8)),
                    7 => std_logic_vector(to_unsigned( 25 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=571 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 80, 8)),
                    1 => std_logic_vector(to_unsigned( 37 , 8)),
                    2 => std_logic_vector(to_unsigned( 100 , 8)),
                    3 => std_logic_vector(to_unsigned( 2 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 93 , 8)),
                    6 => std_logic_vector(to_unsigned( 52 , 8)),
                    7 => std_logic_vector(to_unsigned( 25 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=572 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 122 , 8)),
                    3 => std_logic_vector(to_unsigned( 7 , 8)),
                    4 => std_logic_vector(to_unsigned( 42 , 8)),
                    5 => std_logic_vector(to_unsigned( 47 , 8)),
                    6 => std_logic_vector(to_unsigned( 65 , 8)),
                    7 => std_logic_vector(to_unsigned( 105 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=573 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 71, 8)),
                    1 => std_logic_vector(to_unsigned( 110 , 8)),
                    2 => std_logic_vector(to_unsigned( 52 , 8)),
                    3 => std_logic_vector(to_unsigned( 40 , 8)),
                    4 => std_logic_vector(to_unsigned( 105 , 8)),
                    5 => std_logic_vector(to_unsigned( 61 , 8)),
                    6 => std_logic_vector(to_unsigned( 85 , 8)),
                    7 => std_logic_vector(to_unsigned( 98 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=574 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 71, 8)),
                    1 => std_logic_vector(to_unsigned( 110 , 8)),
                    2 => std_logic_vector(to_unsigned( 52 , 8)),
                    3 => std_logic_vector(to_unsigned( 40 , 8)),
                    4 => std_logic_vector(to_unsigned( 105 , 8)),
                    5 => std_logic_vector(to_unsigned( 61 , 8)),
                    6 => std_logic_vector(to_unsigned( 85 , 8)),
                    7 => std_logic_vector(to_unsigned( 98 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=575 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),
                    1 => std_logic_vector(to_unsigned( 61 , 8)),
                    2 => std_logic_vector(to_unsigned( 30 , 8)),
                    3 => std_logic_vector(to_unsigned( 118 , 8)),
                    4 => std_logic_vector(to_unsigned( 65 , 8)),
                    5 => std_logic_vector(to_unsigned( 47 , 8)),
                    6 => std_logic_vector(to_unsigned( 69 , 8)),
                    7 => std_logic_vector(to_unsigned( 26 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=576 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),
                    1 => std_logic_vector(to_unsigned( 34 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 21 , 8)),
                    6 => std_logic_vector(to_unsigned( 122 , 8)),
                    7 => std_logic_vector(to_unsigned( 14 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=577 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),
                    1 => std_logic_vector(to_unsigned( 34 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 21 , 8)),
                    6 => std_logic_vector(to_unsigned( 122 , 8)),
                    7 => std_logic_vector(to_unsigned( 14 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=578 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 91, 8)),
                    1 => std_logic_vector(to_unsigned( 6 , 8)),
                    2 => std_logic_vector(to_unsigned( 23 , 8)),
                    3 => std_logic_vector(to_unsigned( 95 , 8)),
                    4 => std_logic_vector(to_unsigned( 34 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=579 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 88, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 113 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 21 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=580 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 88, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 113 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 21 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=581 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 82, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 116 , 8)),
                    3 => std_logic_vector(to_unsigned( 12 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 24 , 8)),
                    6 => std_logic_vector(to_unsigned( 112 , 8)),
                    7 => std_logic_vector(to_unsigned( 20 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=582 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 80, 8)),
                    1 => std_logic_vector(to_unsigned( 71 , 8)),
                    2 => std_logic_vector(to_unsigned( 108 , 8)),
                    3 => std_logic_vector(to_unsigned( 17 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 8 , 8)),
                    6 => std_logic_vector(to_unsigned( 46 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=583 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 80, 8)),
                    1 => std_logic_vector(to_unsigned( 71 , 8)),
                    2 => std_logic_vector(to_unsigned( 108 , 8)),
                    3 => std_logic_vector(to_unsigned( 17 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 8 , 8)),
                    6 => std_logic_vector(to_unsigned( 46 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=584 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 7 , 8)),
                    2 => std_logic_vector(to_unsigned( 115 , 8)),
                    3 => std_logic_vector(to_unsigned( 98 , 8)),
                    4 => std_logic_vector(to_unsigned( 82 , 8)),
                    5 => std_logic_vector(to_unsigned( 46 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=585 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),
                    1 => std_logic_vector(to_unsigned( 45 , 8)),
                    2 => std_logic_vector(to_unsigned( 113 , 8)),
                    3 => std_logic_vector(to_unsigned( 15 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 22 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=586 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),
                    1 => std_logic_vector(to_unsigned( 45 , 8)),
                    2 => std_logic_vector(to_unsigned( 113 , 8)),
                    3 => std_logic_vector(to_unsigned( 15 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 22 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=587 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),
                    1 => std_logic_vector(to_unsigned( 62 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 6 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 110 , 8)),
                    7 => std_logic_vector(to_unsigned( 42 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=588 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 70 , 8)),
                    3 => std_logic_vector(to_unsigned( 45 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 23 , 8)),
                    6 => std_logic_vector(to_unsigned( 28 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=589 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 70 , 8)),
                    3 => std_logic_vector(to_unsigned( 45 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 23 , 8)),
                    6 => std_logic_vector(to_unsigned( 28 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=590 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),
                    1 => std_logic_vector(to_unsigned( 2 , 8)),
                    2 => std_logic_vector(to_unsigned( 27 , 8)),
                    3 => std_logic_vector(to_unsigned( 79 , 8)),
                    4 => std_logic_vector(to_unsigned( 101 , 8)),
                    5 => std_logic_vector(to_unsigned( 42 , 8)),
                    6 => std_logic_vector(to_unsigned( 16 , 8)),
                    7 => std_logic_vector(to_unsigned( 121 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=591 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 106, 8)),
                    1 => std_logic_vector(to_unsigned( 77 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 68 , 8)),
                    4 => std_logic_vector(to_unsigned( 52 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 36 , 8)),
                    7 => std_logic_vector(to_unsigned( 122 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=592 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 106, 8)),
                    1 => std_logic_vector(to_unsigned( 77 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 68 , 8)),
                    4 => std_logic_vector(to_unsigned( 52 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 36 , 8)),
                    7 => std_logic_vector(to_unsigned( 122 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=593 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),
                    1 => std_logic_vector(to_unsigned( 111 , 8)),
                    2 => std_logic_vector(to_unsigned( 6 , 8)),
                    3 => std_logic_vector(to_unsigned( 89 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 26 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=594 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 115 , 8)),
                    2 => std_logic_vector(to_unsigned( 97 , 8)),
                    3 => std_logic_vector(to_unsigned( 66 , 8)),
                    4 => std_logic_vector(to_unsigned( 41 , 8)),
                    5 => std_logic_vector(to_unsigned( 75 , 8)),
                    6 => std_logic_vector(to_unsigned( 35 , 8)),
                    7 => std_logic_vector(to_unsigned( 54 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=595 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 115 , 8)),
                    2 => std_logic_vector(to_unsigned( 97 , 8)),
                    3 => std_logic_vector(to_unsigned( 66 , 8)),
                    4 => std_logic_vector(to_unsigned( 41 , 8)),
                    5 => std_logic_vector(to_unsigned( 75 , 8)),
                    6 => std_logic_vector(to_unsigned( 35 , 8)),
                    7 => std_logic_vector(to_unsigned( 54 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=596 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 54 , 8)),
                    2 => std_logic_vector(to_unsigned( 93 , 8)),
                    3 => std_logic_vector(to_unsigned( 44 , 8)),
                    4 => std_logic_vector(to_unsigned( 24 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 16 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=597 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),
                    1 => std_logic_vector(to_unsigned( 63 , 8)),
                    2 => std_logic_vector(to_unsigned( 22 , 8)),
                    3 => std_logic_vector(to_unsigned( 42 , 8)),
                    4 => std_logic_vector(to_unsigned( 116 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 53 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=598 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),
                    1 => std_logic_vector(to_unsigned( 63 , 8)),
                    2 => std_logic_vector(to_unsigned( 22 , 8)),
                    3 => std_logic_vector(to_unsigned( 42 , 8)),
                    4 => std_logic_vector(to_unsigned( 116 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 53 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=599 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 91 , 8)),
                    2 => std_logic_vector(to_unsigned( 14 , 8)),
                    3 => std_logic_vector(to_unsigned( 112 , 8)),
                    4 => std_logic_vector(to_unsigned( 87 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 97 , 8)),
                    7 => std_logic_vector(to_unsigned( 60 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=600 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 103 , 8)),
                    2 => std_logic_vector(to_unsigned( 6 , 8)),
                    3 => std_logic_vector(to_unsigned( 119 , 8)),
                    4 => std_logic_vector(to_unsigned( 22 , 8)),
                    5 => std_logic_vector(to_unsigned( 93 , 8)),
                    6 => std_logic_vector(to_unsigned( 30 , 8)),
                    7 => std_logic_vector(to_unsigned( 16 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=601 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 103 , 8)),
                    2 => std_logic_vector(to_unsigned( 6 , 8)),
                    3 => std_logic_vector(to_unsigned( 119 , 8)),
                    4 => std_logic_vector(to_unsigned( 22 , 8)),
                    5 => std_logic_vector(to_unsigned( 93 , 8)),
                    6 => std_logic_vector(to_unsigned( 30 , 8)),
                    7 => std_logic_vector(to_unsigned( 16 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=602 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 53, 8)),
                    1 => std_logic_vector(to_unsigned( 81 , 8)),
                    2 => std_logic_vector(to_unsigned( 19 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 29 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=603 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 2, 8)),
                    1 => std_logic_vector(to_unsigned( 72 , 8)),
                    2 => std_logic_vector(to_unsigned( 45 , 8)),
                    3 => std_logic_vector(to_unsigned( 84 , 8)),
                    4 => std_logic_vector(to_unsigned( 116 , 8)),
                    5 => std_logic_vector(to_unsigned( 22 , 8)),
                    6 => std_logic_vector(to_unsigned( 105 , 8)),
                    7 => std_logic_vector(to_unsigned( 64 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=604 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 2, 8)),
                    1 => std_logic_vector(to_unsigned( 72 , 8)),
                    2 => std_logic_vector(to_unsigned( 45 , 8)),
                    3 => std_logic_vector(to_unsigned( 84 , 8)),
                    4 => std_logic_vector(to_unsigned( 116 , 8)),
                    5 => std_logic_vector(to_unsigned( 22 , 8)),
                    6 => std_logic_vector(to_unsigned( 105 , 8)),
                    7 => std_logic_vector(to_unsigned( 64 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=605 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 70, 8)),
                    1 => std_logic_vector(to_unsigned( 23 , 8)),
                    2 => std_logic_vector(to_unsigned( 116 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 14 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=606 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 31 , 8)),
                    3 => std_logic_vector(to_unsigned( 65 , 8)),
                    4 => std_logic_vector(to_unsigned( 88 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 54 , 8)),
                    7 => std_logic_vector(to_unsigned( 120 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=607 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 31 , 8)),
                    3 => std_logic_vector(to_unsigned( 65 , 8)),
                    4 => std_logic_vector(to_unsigned( 88 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 54 , 8)),
                    7 => std_logic_vector(to_unsigned( 120 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=608 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 113, 8)),
                    1 => std_logic_vector(to_unsigned( 3 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 57 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 102 , 8)),
                    6 => std_logic_vector(to_unsigned( 18 , 8)),
                    7 => std_logic_vector(to_unsigned( 122 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=609 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),
                    1 => std_logic_vector(to_unsigned( 19 , 8)),
                    2 => std_logic_vector(to_unsigned( 114 , 8)),
                    3 => std_logic_vector(to_unsigned( 12 , 8)),
                    4 => std_logic_vector(to_unsigned( 52 , 8)),
                    5 => std_logic_vector(to_unsigned( 102 , 8)),
                    6 => std_logic_vector(to_unsigned( 68 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=610 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),
                    1 => std_logic_vector(to_unsigned( 19 , 8)),
                    2 => std_logic_vector(to_unsigned( 114 , 8)),
                    3 => std_logic_vector(to_unsigned( 12 , 8)),
                    4 => std_logic_vector(to_unsigned( 52 , 8)),
                    5 => std_logic_vector(to_unsigned( 102 , 8)),
                    6 => std_logic_vector(to_unsigned( 68 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=611 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 105, 8)),
                    1 => std_logic_vector(to_unsigned( 59 , 8)),
                    2 => std_logic_vector(to_unsigned( 28 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 65 , 8)),
                    5 => std_logic_vector(to_unsigned( 10 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 21 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=612 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 62, 8)),
                    1 => std_logic_vector(to_unsigned( 81 , 8)),
                    2 => std_logic_vector(to_unsigned( 122 , 8)),
                    3 => std_logic_vector(to_unsigned( 91 , 8)),
                    4 => std_logic_vector(to_unsigned( 96 , 8)),
                    5 => std_logic_vector(to_unsigned( 30 , 8)),
                    6 => std_logic_vector(to_unsigned( 22 , 8)),
                    7 => std_logic_vector(to_unsigned( 42 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=613 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 62, 8)),
                    1 => std_logic_vector(to_unsigned( 81 , 8)),
                    2 => std_logic_vector(to_unsigned( 122 , 8)),
                    3 => std_logic_vector(to_unsigned( 91 , 8)),
                    4 => std_logic_vector(to_unsigned( 96 , 8)),
                    5 => std_logic_vector(to_unsigned( 30 , 8)),
                    6 => std_logic_vector(to_unsigned( 22 , 8)),
                    7 => std_logic_vector(to_unsigned( 42 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=614 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 121 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 88 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=615 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 27 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 37 , 8)),
                    5 => std_logic_vector(to_unsigned( 33 , 8)),
                    6 => std_logic_vector(to_unsigned( 49 , 8)),
                    7 => std_logic_vector(to_unsigned( 88 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=616 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 27 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 37 , 8)),
                    5 => std_logic_vector(to_unsigned( 33 , 8)),
                    6 => std_logic_vector(to_unsigned( 49 , 8)),
                    7 => std_logic_vector(to_unsigned( 88 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=617 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 37 , 8)),
                    2 => std_logic_vector(to_unsigned( 52 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 108 , 8)),
                    5 => std_logic_vector(to_unsigned( 88 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 65 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=618 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),
                    1 => std_logic_vector(to_unsigned( 16 , 8)),
                    2 => std_logic_vector(to_unsigned( 35 , 8)),
                    3 => std_logic_vector(to_unsigned( 61 , 8)),
                    4 => std_logic_vector(to_unsigned( 11 , 8)),
                    5 => std_logic_vector(to_unsigned( 119 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 112 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=619 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),
                    1 => std_logic_vector(to_unsigned( 16 , 8)),
                    2 => std_logic_vector(to_unsigned( 35 , 8)),
                    3 => std_logic_vector(to_unsigned( 61 , 8)),
                    4 => std_logic_vector(to_unsigned( 11 , 8)),
                    5 => std_logic_vector(to_unsigned( 119 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 112 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=620 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 34 , 8)),
                    2 => std_logic_vector(to_unsigned( 39 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 5 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 14 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=621 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 33 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 76 , 8)),
                    5 => std_logic_vector(to_unsigned( 62 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 118 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=622 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 33 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 76 , 8)),
                    5 => std_logic_vector(to_unsigned( 62 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 118 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=623 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 90, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 6 , 8)),
                    3 => std_logic_vector(to_unsigned( 106 , 8)),
                    4 => std_logic_vector(to_unsigned( 97 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 14 , 8)),
                    7 => std_logic_vector(to_unsigned( 40 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=624 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 21 , 8)),
                    2 => std_logic_vector(to_unsigned( 104 , 8)),
                    3 => std_logic_vector(to_unsigned( 77 , 8)),
                    4 => std_logic_vector(to_unsigned( 119 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 7 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=625 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 21 , 8)),
                    2 => std_logic_vector(to_unsigned( 104 , 8)),
                    3 => std_logic_vector(to_unsigned( 77 , 8)),
                    4 => std_logic_vector(to_unsigned( 119 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 7 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=626 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 81, 8)),
                    1 => std_logic_vector(to_unsigned( 124 , 8)),
                    2 => std_logic_vector(to_unsigned( 91 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 21 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=627 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 82, 8)),
                    1 => std_logic_vector(to_unsigned( 114 , 8)),
                    2 => std_logic_vector(to_unsigned( 101 , 8)),
                    3 => std_logic_vector(to_unsigned( 53 , 8)),
                    4 => std_logic_vector(to_unsigned( 48 , 8)),
                    5 => std_logic_vector(to_unsigned( 39 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=628 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 82, 8)),
                    1 => std_logic_vector(to_unsigned( 114 , 8)),
                    2 => std_logic_vector(to_unsigned( 101 , 8)),
                    3 => std_logic_vector(to_unsigned( 53 , 8)),
                    4 => std_logic_vector(to_unsigned( 48 , 8)),
                    5 => std_logic_vector(to_unsigned( 39 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=629 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 16, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 31 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 37 , 8)),
                    6 => std_logic_vector(to_unsigned( 24 , 8)),
                    7 => std_logic_vector(to_unsigned( 118 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=630 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 40, 8)),
                    1 => std_logic_vector(to_unsigned( 71 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 87 , 8)),
                    5 => std_logic_vector(to_unsigned( 60 , 8)),
                    6 => std_logic_vector(to_unsigned( 24 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=631 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 40, 8)),
                    1 => std_logic_vector(to_unsigned( 71 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 87 , 8)),
                    5 => std_logic_vector(to_unsigned( 60 , 8)),
                    6 => std_logic_vector(to_unsigned( 24 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=632 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 38 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 85 , 8)),
                    5 => std_logic_vector(to_unsigned( 74 , 8)),
                    6 => std_logic_vector(to_unsigned( 124 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=633 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 124 , 8)),
                    2 => std_logic_vector(to_unsigned( 64 , 8)),
                    3 => std_logic_vector(to_unsigned( 55 , 8)),
                    4 => std_logic_vector(to_unsigned( 38 , 8)),
                    5 => std_logic_vector(to_unsigned( 90 , 8)),
                    6 => std_logic_vector(to_unsigned( 109 , 8)),
                    7 => std_logic_vector(to_unsigned( 117 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=634 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 124 , 8)),
                    2 => std_logic_vector(to_unsigned( 64 , 8)),
                    3 => std_logic_vector(to_unsigned( 55 , 8)),
                    4 => std_logic_vector(to_unsigned( 38 , 8)),
                    5 => std_logic_vector(to_unsigned( 90 , 8)),
                    6 => std_logic_vector(to_unsigned( 109 , 8)),
                    7 => std_logic_vector(to_unsigned( 117 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=635 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 47 , 8)),
                    2 => std_logic_vector(to_unsigned( 86 , 8)),
                    3 => std_logic_vector(to_unsigned( 26 , 8)),
                    4 => std_logic_vector(to_unsigned( 114 , 8)),
                    5 => std_logic_vector(to_unsigned( 68 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 107 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=636 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),
                    1 => std_logic_vector(to_unsigned( 119 , 8)),
                    2 => std_logic_vector(to_unsigned( 88 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 28 , 8)),
                    6 => std_logic_vector(to_unsigned( 107 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=637 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),
                    1 => std_logic_vector(to_unsigned( 119 , 8)),
                    2 => std_logic_vector(to_unsigned( 88 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 28 , 8)),
                    6 => std_logic_vector(to_unsigned( 107 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=638 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),
                    1 => std_logic_vector(to_unsigned( 98 , 8)),
                    2 => std_logic_vector(to_unsigned( 30 , 8)),
                    3 => std_logic_vector(to_unsigned( 45 , 8)),
                    4 => std_logic_vector(to_unsigned( 41 , 8)),
                    5 => std_logic_vector(to_unsigned( 19 , 8)),
                    6 => std_logic_vector(to_unsigned( 114 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=639 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 45 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 116 , 8)),
                    5 => std_logic_vector(to_unsigned( 95 , 8)),
                    6 => std_logic_vector(to_unsigned( 107 , 8)),
                    7 => std_logic_vector(to_unsigned( 7 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=640 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 45 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 116 , 8)),
                    5 => std_logic_vector(to_unsigned( 95 , 8)),
                    6 => std_logic_vector(to_unsigned( 107 , 8)),
                    7 => std_logic_vector(to_unsigned( 7 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=641 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 38, 8)),
                    1 => std_logic_vector(to_unsigned( 52 , 8)),
                    2 => std_logic_vector(to_unsigned( 46 , 8)),
                    3 => std_logic_vector(to_unsigned( 84 , 8)),
                    4 => std_logic_vector(to_unsigned( 92 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 27 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=642 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),
                    1 => std_logic_vector(to_unsigned( 79 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 99 , 8)),
                    4 => std_logic_vector(to_unsigned( 64 , 8)),
                    5 => std_logic_vector(to_unsigned( 33 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 115 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=643 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),
                    1 => std_logic_vector(to_unsigned( 79 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 99 , 8)),
                    4 => std_logic_vector(to_unsigned( 64 , 8)),
                    5 => std_logic_vector(to_unsigned( 33 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 115 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=644 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 20, 8)),
                    1 => std_logic_vector(to_unsigned( 108 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 8 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 124 , 8)),
                    7 => std_logic_vector(to_unsigned( 96 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=645 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 5 , 8)),
                    4 => std_logic_vector(to_unsigned( 77 , 8)),
                    5 => std_logic_vector(to_unsigned( 60 , 8)),
                    6 => std_logic_vector(to_unsigned( 113 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=646 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 5 , 8)),
                    4 => std_logic_vector(to_unsigned( 77 , 8)),
                    5 => std_logic_vector(to_unsigned( 60 , 8)),
                    6 => std_logic_vector(to_unsigned( 113 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=647 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 38, 8)),
                    1 => std_logic_vector(to_unsigned( 105 , 8)),
                    2 => std_logic_vector(to_unsigned( 42 , 8)),
                    3 => std_logic_vector(to_unsigned( 118 , 8)),
                    4 => std_logic_vector(to_unsigned( 84 , 8)),
                    5 => std_logic_vector(to_unsigned( 18 , 8)),
                    6 => std_logic_vector(to_unsigned( 76 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=648 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 6 , 8)),
                    2 => std_logic_vector(to_unsigned( 96 , 8)),
                    3 => std_logic_vector(to_unsigned( 16 , 8)),
                    4 => std_logic_vector(to_unsigned( 38 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=649 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 6 , 8)),
                    2 => std_logic_vector(to_unsigned( 96 , 8)),
                    3 => std_logic_vector(to_unsigned( 16 , 8)),
                    4 => std_logic_vector(to_unsigned( 38 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=650 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),
                    1 => std_logic_vector(to_unsigned( 94 , 8)),
                    2 => std_logic_vector(to_unsigned( 85 , 8)),
                    3 => std_logic_vector(to_unsigned( 45 , 8)),
                    4 => std_logic_vector(to_unsigned( 60 , 8)),
                    5 => std_logic_vector(to_unsigned( 22 , 8)),
                    6 => std_logic_vector(to_unsigned( 28 , 8)),
                    7 => std_logic_vector(to_unsigned( 69 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=651 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),
                    1 => std_logic_vector(to_unsigned( 8 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 50 , 8)),
                    6 => std_logic_vector(to_unsigned( 98 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=652 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),
                    1 => std_logic_vector(to_unsigned( 8 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 50 , 8)),
                    6 => std_logic_vector(to_unsigned( 98 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=653 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 46 , 8)),
                    3 => std_logic_vector(to_unsigned( 16 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 66 , 8)),
                    7 => std_logic_vector(to_unsigned( 75 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=654 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),
                    1 => std_logic_vector(to_unsigned( 44 , 8)),
                    2 => std_logic_vector(to_unsigned( 62 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 23 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=655 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),
                    1 => std_logic_vector(to_unsigned( 44 , 8)),
                    2 => std_logic_vector(to_unsigned( 62 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 23 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=656 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 101 , 8)),
                    2 => std_logic_vector(to_unsigned( 53 , 8)),
                    3 => std_logic_vector(to_unsigned( 83 , 8)),
                    4 => std_logic_vector(to_unsigned( 87 , 8)),
                    5 => std_logic_vector(to_unsigned( 34 , 8)),
                    6 => std_logic_vector(to_unsigned( 2 , 8)),
                    7 => std_logic_vector(to_unsigned( 94 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=657 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 112 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 91 , 8)),
                    5 => std_logic_vector(to_unsigned( 102 , 8)),
                    6 => std_logic_vector(to_unsigned( 13 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=658 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 112 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 91 , 8)),
                    5 => std_logic_vector(to_unsigned( 102 , 8)),
                    6 => std_logic_vector(to_unsigned( 13 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=659 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),
                    1 => std_logic_vector(to_unsigned( 80 , 8)),
                    2 => std_logic_vector(to_unsigned( 106 , 8)),
                    3 => std_logic_vector(to_unsigned( 2 , 8)),
                    4 => std_logic_vector(to_unsigned( 120 , 8)),
                    5 => std_logic_vector(to_unsigned( 47 , 8)),
                    6 => std_logic_vector(to_unsigned( 33 , 8)),
                    7 => std_logic_vector(to_unsigned( 75 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=660 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 47, 8)),
                    1 => std_logic_vector(to_unsigned( 107 , 8)),
                    2 => std_logic_vector(to_unsigned( 28 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 24 , 8)),
                    5 => std_logic_vector(to_unsigned( 83 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 58 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=661 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 47, 8)),
                    1 => std_logic_vector(to_unsigned( 107 , 8)),
                    2 => std_logic_vector(to_unsigned( 28 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 24 , 8)),
                    5 => std_logic_vector(to_unsigned( 83 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 58 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=662 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),
                    1 => std_logic_vector(to_unsigned( 89 , 8)),
                    2 => std_logic_vector(to_unsigned( 32 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 6 , 8)),
                    5 => std_logic_vector(to_unsigned( 77 , 8)),
                    6 => std_logic_vector(to_unsigned( 51 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=663 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 61 , 8)),
                    4 => std_logic_vector(to_unsigned( 121 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 19 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=664 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 61 , 8)),
                    4 => std_logic_vector(to_unsigned( 121 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 19 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=665 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),
                    1 => std_logic_vector(to_unsigned( 82 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 8 , 8)),
                    4 => std_logic_vector(to_unsigned( 73 , 8)),
                    5 => std_logic_vector(to_unsigned( 52 , 8)),
                    6 => std_logic_vector(to_unsigned( 87 , 8)),
                    7 => std_logic_vector(to_unsigned( 108 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=666 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 58, 8)),
                    1 => std_logic_vector(to_unsigned( 48 , 8)),
                    2 => std_logic_vector(to_unsigned( 121 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 43 , 8)),
                    5 => std_logic_vector(to_unsigned( 109 , 8)),
                    6 => std_logic_vector(to_unsigned( 87 , 8)),
                    7 => std_logic_vector(to_unsigned( 103 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=667 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 58, 8)),
                    1 => std_logic_vector(to_unsigned( 48 , 8)),
                    2 => std_logic_vector(to_unsigned( 121 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 43 , 8)),
                    5 => std_logic_vector(to_unsigned( 109 , 8)),
                    6 => std_logic_vector(to_unsigned( 87 , 8)),
                    7 => std_logic_vector(to_unsigned( 103 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=668 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 70 , 8)),
                    3 => std_logic_vector(to_unsigned( 119 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 83 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 108 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=669 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 82, 8)),
                    1 => std_logic_vector(to_unsigned( 66 , 8)),
                    2 => std_logic_vector(to_unsigned( 98 , 8)),
                    3 => std_logic_vector(to_unsigned( 121 , 8)),
                    4 => std_logic_vector(to_unsigned( 26 , 8)),
                    5 => std_logic_vector(to_unsigned( 49 , 8)),
                    6 => std_logic_vector(to_unsigned( 21 , 8)),
                    7 => std_logic_vector(to_unsigned( 38 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=670 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 82, 8)),
                    1 => std_logic_vector(to_unsigned( 66 , 8)),
                    2 => std_logic_vector(to_unsigned( 98 , 8)),
                    3 => std_logic_vector(to_unsigned( 121 , 8)),
                    4 => std_logic_vector(to_unsigned( 26 , 8)),
                    5 => std_logic_vector(to_unsigned( 49 , 8)),
                    6 => std_logic_vector(to_unsigned( 21 , 8)),
                    7 => std_logic_vector(to_unsigned( 38 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=671 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 40, 8)),
                    1 => std_logic_vector(to_unsigned( 101 , 8)),
                    2 => std_logic_vector(to_unsigned( 56 , 8)),
                    3 => std_logic_vector(to_unsigned( 116 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 120 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=672 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 50 , 8)),
                    3 => std_logic_vector(to_unsigned( 68 , 8)),
                    4 => std_logic_vector(to_unsigned( 63 , 8)),
                    5 => std_logic_vector(to_unsigned( 42 , 8)),
                    6 => std_logic_vector(to_unsigned( 15 , 8)),
                    7 => std_logic_vector(to_unsigned( 29 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=673 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 50 , 8)),
                    3 => std_logic_vector(to_unsigned( 68 , 8)),
                    4 => std_logic_vector(to_unsigned( 63 , 8)),
                    5 => std_logic_vector(to_unsigned( 42 , 8)),
                    6 => std_logic_vector(to_unsigned( 15 , 8)),
                    7 => std_logic_vector(to_unsigned( 29 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=674 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),
                    1 => std_logic_vector(to_unsigned( 60 , 8)),
                    2 => std_logic_vector(to_unsigned( 1 , 8)),
                    3 => std_logic_vector(to_unsigned( 86 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 72 , 8)),
                    6 => std_logic_vector(to_unsigned( 120 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=675 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 95 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 64 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=676 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 95 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 64 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=677 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 100 , 8)),
                    2 => std_logic_vector(to_unsigned( 40 , 8)),
                    3 => std_logic_vector(to_unsigned( 119 , 8)),
                    4 => std_logic_vector(to_unsigned( 82 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 63 , 8)),
                    7 => std_logic_vector(to_unsigned( 112 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=678 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 105, 8)),
                    1 => std_logic_vector(to_unsigned( 44 , 8)),
                    2 => std_logic_vector(to_unsigned( 53 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 6 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 123 , 8)),
                    7 => std_logic_vector(to_unsigned( 26 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=679 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 105, 8)),
                    1 => std_logic_vector(to_unsigned( 44 , 8)),
                    2 => std_logic_vector(to_unsigned( 53 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 6 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 123 , 8)),
                    7 => std_logic_vector(to_unsigned( 26 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=680 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 116 , 8)),
                    3 => std_logic_vector(to_unsigned( 124 , 8)),
                    4 => std_logic_vector(to_unsigned( 17 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 25 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=681 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 54 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 23 , 8)),
                    5 => std_logic_vector(to_unsigned( 46 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=682 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 54 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 23 , 8)),
                    5 => std_logic_vector(to_unsigned( 46 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=683 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 72, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 93 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 101 , 8)),
                    5 => std_logic_vector(to_unsigned( 14 , 8)),
                    6 => std_logic_vector(to_unsigned( 116 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=684 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 99, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 106 , 8)),
                    4 => std_logic_vector(to_unsigned( 92 , 8)),
                    5 => std_logic_vector(to_unsigned( 22 , 8)),
                    6 => std_logic_vector(to_unsigned( 49 , 8)),
                    7 => std_logic_vector(to_unsigned( 59 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=685 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 99, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 106 , 8)),
                    4 => std_logic_vector(to_unsigned( 92 , 8)),
                    5 => std_logic_vector(to_unsigned( 22 , 8)),
                    6 => std_logic_vector(to_unsigned( 49 , 8)),
                    7 => std_logic_vector(to_unsigned( 59 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=686 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),
                    1 => std_logic_vector(to_unsigned( 53 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 111 , 8)),
                    6 => std_logic_vector(to_unsigned( 115 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=687 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 20, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 111 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 3 , 8)),
                    5 => std_logic_vector(to_unsigned( 28 , 8)),
                    6 => std_logic_vector(to_unsigned( 92 , 8)),
                    7 => std_logic_vector(to_unsigned( 78 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=688 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 20, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 111 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 3 , 8)),
                    5 => std_logic_vector(to_unsigned( 28 , 8)),
                    6 => std_logic_vector(to_unsigned( 92 , 8)),
                    7 => std_logic_vector(to_unsigned( 78 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=689 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 5 , 8)),
                    2 => std_logic_vector(to_unsigned( 93 , 8)),
                    3 => std_logic_vector(to_unsigned( 113 , 8)),
                    4 => std_logic_vector(to_unsigned( 47 , 8)),
                    5 => std_logic_vector(to_unsigned( 38 , 8)),
                    6 => std_logic_vector(to_unsigned( 61 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=690 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 27 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 57 , 8)),
                    4 => std_logic_vector(to_unsigned( 63 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=691 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 27 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 57 , 8)),
                    4 => std_logic_vector(to_unsigned( 63 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=692 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 73, 8)),
                    1 => std_logic_vector(to_unsigned( 123 , 8)),
                    2 => std_logic_vector(to_unsigned( 28 , 8)),
                    3 => std_logic_vector(to_unsigned( 81 , 8)),
                    4 => std_logic_vector(to_unsigned( 119 , 8)),
                    5 => std_logic_vector(to_unsigned( 91 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 99 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=693 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 83, 8)),
                    1 => std_logic_vector(to_unsigned( 104 , 8)),
                    2 => std_logic_vector(to_unsigned( 120 , 8)),
                    3 => std_logic_vector(to_unsigned( 97 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 54 , 8)),
                    7 => std_logic_vector(to_unsigned( 71 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=694 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 83, 8)),
                    1 => std_logic_vector(to_unsigned( 104 , 8)),
                    2 => std_logic_vector(to_unsigned( 120 , 8)),
                    3 => std_logic_vector(to_unsigned( 97 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 54 , 8)),
                    7 => std_logic_vector(to_unsigned( 71 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=695 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 109, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 70 , 8)),
                    3 => std_logic_vector(to_unsigned( 20 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 50 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=696 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 80, 8)),
                    1 => std_logic_vector(to_unsigned( 25 , 8)),
                    2 => std_logic_vector(to_unsigned( 57 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 112 , 8)),
                    6 => std_logic_vector(to_unsigned( 13 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=697 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 80, 8)),
                    1 => std_logic_vector(to_unsigned( 25 , 8)),
                    2 => std_logic_vector(to_unsigned( 57 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 112 , 8)),
                    6 => std_logic_vector(to_unsigned( 13 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=698 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),
                    1 => std_logic_vector(to_unsigned( 94 , 8)),
                    2 => std_logic_vector(to_unsigned( 38 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 114 , 8)),
                    5 => std_logic_vector(to_unsigned( 14 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 122 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=699 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 61 , 8)),
                    2 => std_logic_vector(to_unsigned( 21 , 8)),
                    3 => std_logic_vector(to_unsigned( 97 , 8)),
                    4 => std_logic_vector(to_unsigned( 47 , 8)),
                    5 => std_logic_vector(to_unsigned( 115 , 8)),
                    6 => std_logic_vector(to_unsigned( 41 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=700 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 61 , 8)),
                    2 => std_logic_vector(to_unsigned( 21 , 8)),
                    3 => std_logic_vector(to_unsigned( 97 , 8)),
                    4 => std_logic_vector(to_unsigned( 47 , 8)),
                    5 => std_logic_vector(to_unsigned( 115 , 8)),
                    6 => std_logic_vector(to_unsigned( 41 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=701 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 122 , 8)),
                    3 => std_logic_vector(to_unsigned( 28 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 22 , 8)),
                    6 => std_logic_vector(to_unsigned( 67 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=702 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),
                    1 => std_logic_vector(to_unsigned( 94 , 8)),
                    2 => std_logic_vector(to_unsigned( 10 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 72 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 27 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=703 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),
                    1 => std_logic_vector(to_unsigned( 94 , 8)),
                    2 => std_logic_vector(to_unsigned( 10 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 72 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 27 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=704 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),
                    1 => std_logic_vector(to_unsigned( 60 , 8)),
                    2 => std_logic_vector(to_unsigned( 109 , 8)),
                    3 => std_logic_vector(to_unsigned( 122 , 8)),
                    4 => std_logic_vector(to_unsigned( 2 , 8)),
                    5 => std_logic_vector(to_unsigned( 84 , 8)),
                    6 => std_logic_vector(to_unsigned( 12 , 8)),
                    7 => std_logic_vector(to_unsigned( 70 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=705 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),
                    1 => std_logic_vector(to_unsigned( 117 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 65 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 92 , 8)),
                    7 => std_logic_vector(to_unsigned( 46 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=706 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),
                    1 => std_logic_vector(to_unsigned( 117 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 65 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 92 , 8)),
                    7 => std_logic_vector(to_unsigned( 46 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=707 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 27 , 8)),
                    2 => std_logic_vector(to_unsigned( 75 , 8)),
                    3 => std_logic_vector(to_unsigned( 120 , 8)),
                    4 => std_logic_vector(to_unsigned( 59 , 8)),
                    5 => std_logic_vector(to_unsigned( 11 , 8)),
                    6 => std_logic_vector(to_unsigned( 32 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=708 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 81, 8)),
                    1 => std_logic_vector(to_unsigned( 31 , 8)),
                    2 => std_logic_vector(to_unsigned( 97 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 124 , 8)),
                    5 => std_logic_vector(to_unsigned( 17 , 8)),
                    6 => std_logic_vector(to_unsigned( 48 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=709 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 81, 8)),
                    1 => std_logic_vector(to_unsigned( 31 , 8)),
                    2 => std_logic_vector(to_unsigned( 97 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 124 , 8)),
                    5 => std_logic_vector(to_unsigned( 17 , 8)),
                    6 => std_logic_vector(to_unsigned( 48 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=710 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 32 , 8)),
                    3 => std_logic_vector(to_unsigned( 59 , 8)),
                    4 => std_logic_vector(to_unsigned( 118 , 8)),
                    5 => std_logic_vector(to_unsigned( 123 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=711 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 91, 8)),
                    1 => std_logic_vector(to_unsigned( 70 , 8)),
                    2 => std_logic_vector(to_unsigned( 50 , 8)),
                    3 => std_logic_vector(to_unsigned( 21 , 8)),
                    4 => std_logic_vector(to_unsigned( 114 , 8)),
                    5 => std_logic_vector(to_unsigned( 118 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 27 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=712 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 91, 8)),
                    1 => std_logic_vector(to_unsigned( 70 , 8)),
                    2 => std_logic_vector(to_unsigned( 50 , 8)),
                    3 => std_logic_vector(to_unsigned( 21 , 8)),
                    4 => std_logic_vector(to_unsigned( 114 , 8)),
                    5 => std_logic_vector(to_unsigned( 118 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 27 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=713 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 16, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 34 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 94 , 8)),
                    5 => std_logic_vector(to_unsigned( 102 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 82 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=714 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 45, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 76 , 8)),
                    5 => std_logic_vector(to_unsigned( 33 , 8)),
                    6 => std_logic_vector(to_unsigned( 16 , 8)),
                    7 => std_logic_vector(to_unsigned( 117 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=715 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 45, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 76 , 8)),
                    5 => std_logic_vector(to_unsigned( 33 , 8)),
                    6 => std_logic_vector(to_unsigned( 16 , 8)),
                    7 => std_logic_vector(to_unsigned( 117 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=716 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 62, 8)),
                    1 => std_logic_vector(to_unsigned( 82 , 8)),
                    2 => std_logic_vector(to_unsigned( 50 , 8)),
                    3 => std_logic_vector(to_unsigned( 109 , 8)),
                    4 => std_logic_vector(to_unsigned( 119 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=717 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),
                    1 => std_logic_vector(to_unsigned( 68 , 8)),
                    2 => std_logic_vector(to_unsigned( 80 , 8)),
                    3 => std_logic_vector(to_unsigned( 46 , 8)),
                    4 => std_logic_vector(to_unsigned( 6 , 8)),
                    5 => std_logic_vector(to_unsigned( 41 , 8)),
                    6 => std_logic_vector(to_unsigned( 18 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=718 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),
                    1 => std_logic_vector(to_unsigned( 68 , 8)),
                    2 => std_logic_vector(to_unsigned( 80 , 8)),
                    3 => std_logic_vector(to_unsigned( 46 , 8)),
                    4 => std_logic_vector(to_unsigned( 6 , 8)),
                    5 => std_logic_vector(to_unsigned( 41 , 8)),
                    6 => std_logic_vector(to_unsigned( 18 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=719 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),
                    1 => std_logic_vector(to_unsigned( 61 , 8)),
                    2 => std_logic_vector(to_unsigned( 67 , 8)),
                    3 => std_logic_vector(to_unsigned( 39 , 8)),
                    4 => std_logic_vector(to_unsigned( 75 , 8)),
                    5 => std_logic_vector(to_unsigned( 99 , 8)),
                    6 => std_logic_vector(to_unsigned( 4 , 8)),
                    7 => std_logic_vector(to_unsigned( 25 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=720 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 93 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 87 , 8)),
                    5 => std_logic_vector(to_unsigned( 110 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 116 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=721 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 93 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 87 , 8)),
                    5 => std_logic_vector(to_unsigned( 110 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 116 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=722 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 109, 8)),
                    1 => std_logic_vector(to_unsigned( 53 , 8)),
                    2 => std_logic_vector(to_unsigned( 88 , 8)),
                    3 => std_logic_vector(to_unsigned( 12 , 8)),
                    4 => std_logic_vector(to_unsigned( 41 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 28 , 8)),
                    7 => std_logic_vector(to_unsigned( 100 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=723 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 75 , 8)),
                    2 => std_logic_vector(to_unsigned( 21 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 108 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 79 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=724 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 75 , 8)),
                    2 => std_logic_vector(to_unsigned( 21 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 108 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 79 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=725 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 76, 8)),
                    1 => std_logic_vector(to_unsigned( 30 , 8)),
                    2 => std_logic_vector(to_unsigned( 57 , 8)),
                    3 => std_logic_vector(to_unsigned( 46 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 88 , 8)),
                    7 => std_logic_vector(to_unsigned( 36 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=726 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 73 , 8)),
                    3 => std_logic_vector(to_unsigned( 107 , 8)),
                    4 => std_logic_vector(to_unsigned( 12 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 5 , 8)),
                    7 => std_logic_vector(to_unsigned( 31 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=727 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 73 , 8)),
                    3 => std_logic_vector(to_unsigned( 107 , 8)),
                    4 => std_logic_vector(to_unsigned( 12 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 5 , 8)),
                    7 => std_logic_vector(to_unsigned( 31 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=728 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 84 , 8)),
                    2 => std_logic_vector(to_unsigned( 22 , 8)),
                    3 => std_logic_vector(to_unsigned( 43 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 8 , 8)),
                    6 => std_logic_vector(to_unsigned( 92 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=729 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 41 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=730 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 41 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=731 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 63 , 8)),
                    2 => std_logic_vector(to_unsigned( 3 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 57 , 8)),
                    5 => std_logic_vector(to_unsigned( 112 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 10 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=732 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 14 , 8)),
                    2 => std_logic_vector(to_unsigned( 63 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 4 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 102 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=733 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 14 , 8)),
                    2 => std_logic_vector(to_unsigned( 63 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 4 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 102 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=734 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 99, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 56 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 3 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 38 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=735 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 52 , 8)),
                    3 => std_logic_vector(to_unsigned( 114 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 48 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=736 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 52 , 8)),
                    3 => std_logic_vector(to_unsigned( 114 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 48 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=737 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),
                    1 => std_logic_vector(to_unsigned( 94 , 8)),
                    2 => std_logic_vector(to_unsigned( 45 , 8)),
                    3 => std_logic_vector(to_unsigned( 23 , 8)),
                    4 => std_logic_vector(to_unsigned( 78 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 1 , 8)),
                    7 => std_logic_vector(to_unsigned( 13 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=738 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 41, 8)),
                    1 => std_logic_vector(to_unsigned( 61 , 8)),
                    2 => std_logic_vector(to_unsigned( 74 , 8)),
                    3 => std_logic_vector(to_unsigned( 5 , 8)),
                    4 => std_logic_vector(to_unsigned( 120 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 104 , 8)),
                    7 => std_logic_vector(to_unsigned( 1 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=739 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 41, 8)),
                    1 => std_logic_vector(to_unsigned( 61 , 8)),
                    2 => std_logic_vector(to_unsigned( 74 , 8)),
                    3 => std_logic_vector(to_unsigned( 5 , 8)),
                    4 => std_logic_vector(to_unsigned( 120 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 104 , 8)),
                    7 => std_logic_vector(to_unsigned( 1 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=740 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),
                    1 => std_logic_vector(to_unsigned( 104 , 8)),
                    2 => std_logic_vector(to_unsigned( 18 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 8 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 87 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=741 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 53, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 48 , 8)),
                    3 => std_logic_vector(to_unsigned( 112 , 8)),
                    4 => std_logic_vector(to_unsigned( 120 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 100 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=742 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 53, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 48 , 8)),
                    3 => std_logic_vector(to_unsigned( 112 , 8)),
                    4 => std_logic_vector(to_unsigned( 120 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 100 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=743 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 90 , 8)),
                    3 => std_logic_vector(to_unsigned( 49 , 8)),
                    4 => std_logic_vector(to_unsigned( 7 , 8)),
                    5 => std_logic_vector(to_unsigned( 117 , 8)),
                    6 => std_logic_vector(to_unsigned( 105 , 8)),
                    7 => std_logic_vector(to_unsigned( 83 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=744 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),
                    1 => std_logic_vector(to_unsigned( 58 , 8)),
                    2 => std_logic_vector(to_unsigned( 69 , 8)),
                    3 => std_logic_vector(to_unsigned( 26 , 8)),
                    4 => std_logic_vector(to_unsigned( 30 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 20 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=745 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),
                    1 => std_logic_vector(to_unsigned( 58 , 8)),
                    2 => std_logic_vector(to_unsigned( 69 , 8)),
                    3 => std_logic_vector(to_unsigned( 26 , 8)),
                    4 => std_logic_vector(to_unsigned( 30 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 20 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=746 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 67, 8)),
                    1 => std_logic_vector(to_unsigned( 21 , 8)),
                    2 => std_logic_vector(to_unsigned( 122 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 82 , 8)),
                    5 => std_logic_vector(to_unsigned( 8 , 8)),
                    6 => std_logic_vector(to_unsigned( 111 , 8)),
                    7 => std_logic_vector(to_unsigned( 104 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=747 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),
                    1 => std_logic_vector(to_unsigned( 71 , 8)),
                    2 => std_logic_vector(to_unsigned( 14 , 8)),
                    3 => std_logic_vector(to_unsigned( 62 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 24 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 36 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=748 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),
                    1 => std_logic_vector(to_unsigned( 71 , 8)),
                    2 => std_logic_vector(to_unsigned( 14 , 8)),
                    3 => std_logic_vector(to_unsigned( 62 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 24 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 36 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=749 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),
                    1 => std_logic_vector(to_unsigned( 53 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 46 , 8)),
                    4 => std_logic_vector(to_unsigned( 6 , 8)),
                    5 => std_logic_vector(to_unsigned( 33 , 8)),
                    6 => std_logic_vector(to_unsigned( 68 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=750 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 80 , 8)),
                    2 => std_logic_vector(to_unsigned( 19 , 8)),
                    3 => std_logic_vector(to_unsigned( 11 , 8)),
                    4 => std_logic_vector(to_unsigned( 51 , 8)),
                    5 => std_logic_vector(to_unsigned( 36 , 8)),
                    6 => std_logic_vector(to_unsigned( 120 , 8)),
                    7 => std_logic_vector(to_unsigned( 62 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=751 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 80 , 8)),
                    2 => std_logic_vector(to_unsigned( 19 , 8)),
                    3 => std_logic_vector(to_unsigned( 11 , 8)),
                    4 => std_logic_vector(to_unsigned( 51 , 8)),
                    5 => std_logic_vector(to_unsigned( 36 , 8)),
                    6 => std_logic_vector(to_unsigned( 120 , 8)),
                    7 => std_logic_vector(to_unsigned( 62 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=752 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 12 , 8)),
                    2 => std_logic_vector(to_unsigned( 83 , 8)),
                    3 => std_logic_vector(to_unsigned( 5 , 8)),
                    4 => std_logic_vector(to_unsigned( 59 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 45 , 8)),
                    7 => std_logic_vector(to_unsigned( 112 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=753 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),
                    1 => std_logic_vector(to_unsigned( 112 , 8)),
                    2 => std_logic_vector(to_unsigned( 91 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 45 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 57 , 8)),
                    7 => std_logic_vector(to_unsigned( 82 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=754 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),
                    1 => std_logic_vector(to_unsigned( 112 , 8)),
                    2 => std_logic_vector(to_unsigned( 91 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 45 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 57 , 8)),
                    7 => std_logic_vector(to_unsigned( 82 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=755 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 17 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 122 , 8)),
                    7 => std_logic_vector(to_unsigned( 81 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=756 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),
                    1 => std_logic_vector(to_unsigned( 29 , 8)),
                    2 => std_logic_vector(to_unsigned( 1 , 8)),
                    3 => std_logic_vector(to_unsigned( 106 , 8)),
                    4 => std_logic_vector(to_unsigned( 72 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=757 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),
                    1 => std_logic_vector(to_unsigned( 29 , 8)),
                    2 => std_logic_vector(to_unsigned( 1 , 8)),
                    3 => std_logic_vector(to_unsigned( 106 , 8)),
                    4 => std_logic_vector(to_unsigned( 72 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=758 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 109, 8)),
                    1 => std_logic_vector(to_unsigned( 18 , 8)),
                    2 => std_logic_vector(to_unsigned( 32 , 8)),
                    3 => std_logic_vector(to_unsigned( 7 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 45 , 8)),
                    7 => std_logic_vector(to_unsigned( 57 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=759 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 58, 8)),
                    1 => std_logic_vector(to_unsigned( 19 , 8)),
                    2 => std_logic_vector(to_unsigned( 70 , 8)),
                    3 => std_logic_vector(to_unsigned( 36 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 26 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=760 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 58, 8)),
                    1 => std_logic_vector(to_unsigned( 19 , 8)),
                    2 => std_logic_vector(to_unsigned( 70 , 8)),
                    3 => std_logic_vector(to_unsigned( 36 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 26 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=761 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 17, 8)),
                    1 => std_logic_vector(to_unsigned( 71 , 8)),
                    2 => std_logic_vector(to_unsigned( 22 , 8)),
                    3 => std_logic_vector(to_unsigned( 76 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 92 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 83 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=762 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),
                    1 => std_logic_vector(to_unsigned( 29 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 123 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 24 , 8)),
                    6 => std_logic_vector(to_unsigned( 60 , 8)),
                    7 => std_logic_vector(to_unsigned( 68 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=763 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),
                    1 => std_logic_vector(to_unsigned( 29 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 123 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 24 , 8)),
                    6 => std_logic_vector(to_unsigned( 60 , 8)),
                    7 => std_logic_vector(to_unsigned( 68 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=764 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 58, 8)),
                    1 => std_logic_vector(to_unsigned( 120 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 25 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 34 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 18 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=765 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 25 , 8)),
                    2 => std_logic_vector(to_unsigned( 106 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 60 , 8)),
                    5 => std_logic_vector(to_unsigned( 54 , 8)),
                    6 => std_logic_vector(to_unsigned( 78 , 8)),
                    7 => std_logic_vector(to_unsigned( 9 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=766 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 25 , 8)),
                    2 => std_logic_vector(to_unsigned( 106 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 60 , 8)),
                    5 => std_logic_vector(to_unsigned( 54 , 8)),
                    6 => std_logic_vector(to_unsigned( 78 , 8)),
                    7 => std_logic_vector(to_unsigned( 9 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=767 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 118 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 98 , 8)),
                    4 => std_logic_vector(to_unsigned( 108 , 8)),
                    5 => std_logic_vector(to_unsigned( 13 , 8)),
                    6 => std_logic_vector(to_unsigned( 102 , 8)),
                    7 => std_logic_vector(to_unsigned( 5 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=768 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 99 , 8)),
                    4 => std_logic_vector(to_unsigned( 123 , 8)),
                    5 => std_logic_vector(to_unsigned( 90 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=769 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 99 , 8)),
                    4 => std_logic_vector(to_unsigned( 123 , 8)),
                    5 => std_logic_vector(to_unsigned( 90 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=770 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),
                    1 => std_logic_vector(to_unsigned( 86 , 8)),
                    2 => std_logic_vector(to_unsigned( 22 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 50 , 8)),
                    6 => std_logic_vector(to_unsigned( 124 , 8)),
                    7 => std_logic_vector(to_unsigned( 56 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=771 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 121 , 8)),
                    4 => std_logic_vector(to_unsigned( 56 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 116 , 8)),
                    7 => std_logic_vector(to_unsigned( 42 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=772 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 121 , 8)),
                    4 => std_logic_vector(to_unsigned( 56 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 116 , 8)),
                    7 => std_logic_vector(to_unsigned( 42 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=773 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 38 , 8)),
                    3 => std_logic_vector(to_unsigned( 3 , 8)),
                    4 => std_logic_vector(to_unsigned( 44 , 8)),
                    5 => std_logic_vector(to_unsigned( 93 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 58 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=774 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 85 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 69 , 8)),
                    5 => std_logic_vector(to_unsigned( 105 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 79 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=775 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 85 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 69 , 8)),
                    5 => std_logic_vector(to_unsigned( 105 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 79 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=776 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 40, 8)),
                    1 => std_logic_vector(to_unsigned( 77 , 8)),
                    2 => std_logic_vector(to_unsigned( 96 , 8)),
                    3 => std_logic_vector(to_unsigned( 29 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 19 , 8)),
                    6 => std_logic_vector(to_unsigned( 50 , 8)),
                    7 => std_logic_vector(to_unsigned( 70 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=777 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),
                    1 => std_logic_vector(to_unsigned( 3 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 121 , 8)),
                    4 => std_logic_vector(to_unsigned( 47 , 8)),
                    5 => std_logic_vector(to_unsigned( 72 , 8)),
                    6 => std_logic_vector(to_unsigned( 67 , 8)),
                    7 => std_logic_vector(to_unsigned( 35 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=778 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),
                    1 => std_logic_vector(to_unsigned( 3 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 121 , 8)),
                    4 => std_logic_vector(to_unsigned( 47 , 8)),
                    5 => std_logic_vector(to_unsigned( 72 , 8)),
                    6 => std_logic_vector(to_unsigned( 67 , 8)),
                    7 => std_logic_vector(to_unsigned( 35 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=779 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 63, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 33 , 8)),
                    3 => std_logic_vector(to_unsigned( 107 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 82 , 8)),
                    6 => std_logic_vector(to_unsigned( 5 , 8)),
                    7 => std_logic_vector(to_unsigned( 87 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=780 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 98 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 103 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 43 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=781 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 98 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 103 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 43 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=782 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 92 , 8)),
                    2 => std_logic_vector(to_unsigned( 46 , 8)),
                    3 => std_logic_vector(to_unsigned( 10 , 8)),
                    4 => std_logic_vector(to_unsigned( 20 , 8)),
                    5 => std_logic_vector(to_unsigned( 122 , 8)),
                    6 => std_logic_vector(to_unsigned( 27 , 8)),
                    7 => std_logic_vector(to_unsigned( 88 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=783 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 78 , 8)),
                    3 => std_logic_vector(to_unsigned( 123 , 8)),
                    4 => std_logic_vector(to_unsigned( 38 , 8)),
                    5 => std_logic_vector(to_unsigned( 5 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 29 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=784 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 78 , 8)),
                    3 => std_logic_vector(to_unsigned( 123 , 8)),
                    4 => std_logic_vector(to_unsigned( 38 , 8)),
                    5 => std_logic_vector(to_unsigned( 5 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 29 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=785 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 76, 8)),
                    1 => std_logic_vector(to_unsigned( 7 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 113 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 62 , 8)),
                    6 => std_logic_vector(to_unsigned( 48 , 8)),
                    7 => std_logic_vector(to_unsigned( 55 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=786 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),
                    1 => std_logic_vector(to_unsigned( 91 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 105 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 35 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=787 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),
                    1 => std_logic_vector(to_unsigned( 91 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 105 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 35 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=788 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 46, 8)),
                    1 => std_logic_vector(to_unsigned( 100 , 8)),
                    2 => std_logic_vector(to_unsigned( 14 , 8)),
                    3 => std_logic_vector(to_unsigned( 8 , 8)),
                    4 => std_logic_vector(to_unsigned( 121 , 8)),
                    5 => std_logic_vector(to_unsigned( 95 , 8)),
                    6 => std_logic_vector(to_unsigned( 59 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=789 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 39 , 8)),
                    3 => std_logic_vector(to_unsigned( 60 , 8)),
                    4 => std_logic_vector(to_unsigned( 84 , 8)),
                    5 => std_logic_vector(to_unsigned( 51 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 105 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=790 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 39 , 8)),
                    3 => std_logic_vector(to_unsigned( 60 , 8)),
                    4 => std_logic_vector(to_unsigned( 84 , 8)),
                    5 => std_logic_vector(to_unsigned( 51 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 105 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=791 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 15 , 8)),
                    4 => std_logic_vector(to_unsigned( 59 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 27 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=792 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 101 , 8)),
                    3 => std_logic_vector(to_unsigned( 65 , 8)),
                    4 => std_logic_vector(to_unsigned( 39 , 8)),
                    5 => std_logic_vector(to_unsigned( 50 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 15 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=793 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 101 , 8)),
                    3 => std_logic_vector(to_unsigned( 65 , 8)),
                    4 => std_logic_vector(to_unsigned( 39 , 8)),
                    5 => std_logic_vector(to_unsigned( 50 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 15 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=794 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),
                    1 => std_logic_vector(to_unsigned( 2 , 8)),
                    2 => std_logic_vector(to_unsigned( 79 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 9 , 8)),
                    5 => std_logic_vector(to_unsigned( 102 , 8)),
                    6 => std_logic_vector(to_unsigned( 29 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=795 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),
                    1 => std_logic_vector(to_unsigned( 63 , 8)),
                    2 => std_logic_vector(to_unsigned( 31 , 8)),
                    3 => std_logic_vector(to_unsigned( 25 , 8)),
                    4 => std_logic_vector(to_unsigned( 73 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 92 , 8)),
                    7 => std_logic_vector(to_unsigned( 18 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=796 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),
                    1 => std_logic_vector(to_unsigned( 63 , 8)),
                    2 => std_logic_vector(to_unsigned( 31 , 8)),
                    3 => std_logic_vector(to_unsigned( 25 , 8)),
                    4 => std_logic_vector(to_unsigned( 73 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 92 , 8)),
                    7 => std_logic_vector(to_unsigned( 18 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=797 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 113, 8)),
                    1 => std_logic_vector(to_unsigned( 121 , 8)),
                    2 => std_logic_vector(to_unsigned( 47 , 8)),
                    3 => std_logic_vector(to_unsigned( 58 , 8)),
                    4 => std_logic_vector(to_unsigned( 24 , 8)),
                    5 => std_logic_vector(to_unsigned( 102 , 8)),
                    6 => std_logic_vector(to_unsigned( 30 , 8)),
                    7 => std_logic_vector(to_unsigned( 4 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=798 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),
                    1 => std_logic_vector(to_unsigned( 31 , 8)),
                    2 => std_logic_vector(to_unsigned( 105 , 8)),
                    3 => std_logic_vector(to_unsigned( 67 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 14 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=799 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),
                    1 => std_logic_vector(to_unsigned( 31 , 8)),
                    2 => std_logic_vector(to_unsigned( 105 , 8)),
                    3 => std_logic_vector(to_unsigned( 67 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 14 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=800 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 46 , 8)),
                    2 => std_logic_vector(to_unsigned( 89 , 8)),
                    3 => std_logic_vector(to_unsigned( 106 , 8)),
                    4 => std_logic_vector(to_unsigned( 101 , 8)),
                    5 => std_logic_vector(to_unsigned( 6 , 8)),
                    6 => std_logic_vector(to_unsigned( 60 , 8)),
                    7 => std_logic_vector(to_unsigned( 24 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=801 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 110, 8)),
                    1 => std_logic_vector(to_unsigned( 16 , 8)),
                    2 => std_logic_vector(to_unsigned( 81 , 8)),
                    3 => std_logic_vector(to_unsigned( 120 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 114 , 8)),
                    7 => std_logic_vector(to_unsigned( 68 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=802 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 110, 8)),
                    1 => std_logic_vector(to_unsigned( 16 , 8)),
                    2 => std_logic_vector(to_unsigned( 81 , 8)),
                    3 => std_logic_vector(to_unsigned( 120 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 114 , 8)),
                    7 => std_logic_vector(to_unsigned( 68 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=803 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),
                    1 => std_logic_vector(to_unsigned( 39 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 75 , 8)),
                    4 => std_logic_vector(to_unsigned( 4 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 59 , 8)),
                    7 => std_logic_vector(to_unsigned( 53 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=804 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 47, 8)),
                    1 => std_logic_vector(to_unsigned( 109 , 8)),
                    2 => std_logic_vector(to_unsigned( 93 , 8)),
                    3 => std_logic_vector(to_unsigned( 23 , 8)),
                    4 => std_logic_vector(to_unsigned( 56 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 88 , 8)),
                    7 => std_logic_vector(to_unsigned( 83 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=805 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 47, 8)),
                    1 => std_logic_vector(to_unsigned( 109 , 8)),
                    2 => std_logic_vector(to_unsigned( 93 , 8)),
                    3 => std_logic_vector(to_unsigned( 23 , 8)),
                    4 => std_logic_vector(to_unsigned( 56 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 88 , 8)),
                    7 => std_logic_vector(to_unsigned( 83 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=806 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 8 , 8)),
                    2 => std_logic_vector(to_unsigned( 68 , 8)),
                    3 => std_logic_vector(to_unsigned( 12 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 78 , 8)),
                    6 => std_logic_vector(to_unsigned( 43 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=807 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 83, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 96 , 8)),
                    4 => std_logic_vector(to_unsigned( 66 , 8)),
                    5 => std_logic_vector(to_unsigned( 88 , 8)),
                    6 => std_logic_vector(to_unsigned( 36 , 8)),
                    7 => std_logic_vector(to_unsigned( 21 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=808 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 83, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 96 , 8)),
                    4 => std_logic_vector(to_unsigned( 66 , 8)),
                    5 => std_logic_vector(to_unsigned( 88 , 8)),
                    6 => std_logic_vector(to_unsigned( 36 , 8)),
                    7 => std_logic_vector(to_unsigned( 21 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=809 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 57 , 8)),
                    2 => std_logic_vector(to_unsigned( 9 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 42 , 8)),
                    5 => std_logic_vector(to_unsigned( 73 , 8)),
                    6 => std_logic_vector(to_unsigned( 87 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=810 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 115 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 37 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 70 , 8)),
                    7 => std_logic_vector(to_unsigned( 28 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=811 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 115 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 37 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 70 , 8)),
                    7 => std_logic_vector(to_unsigned( 28 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=812 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 25, 8)),
                    1 => std_logic_vector(to_unsigned( 84 , 8)),
                    2 => std_logic_vector(to_unsigned( 120 , 8)),
                    3 => std_logic_vector(to_unsigned( 37 , 8)),
                    4 => std_logic_vector(to_unsigned( 19 , 8)),
                    5 => std_logic_vector(to_unsigned( 55 , 8)),
                    6 => std_logic_vector(to_unsigned( 49 , 8)),
                    7 => std_logic_vector(to_unsigned( 62 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=813 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 91 , 8)),
                    2 => std_logic_vector(to_unsigned( 49 , 8)),
                    3 => std_logic_vector(to_unsigned( 116 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 15 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 36 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=814 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 91 , 8)),
                    2 => std_logic_vector(to_unsigned( 49 , 8)),
                    3 => std_logic_vector(to_unsigned( 116 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 15 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 36 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=815 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),
                    1 => std_logic_vector(to_unsigned( 15 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 39 , 8)),
                    5 => std_logic_vector(to_unsigned( 115 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 51 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=816 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),
                    1 => std_logic_vector(to_unsigned( 51 , 8)),
                    2 => std_logic_vector(to_unsigned( 73 , 8)),
                    3 => std_logic_vector(to_unsigned( 20 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 112 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=817 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),
                    1 => std_logic_vector(to_unsigned( 51 , 8)),
                    2 => std_logic_vector(to_unsigned( 73 , 8)),
                    3 => std_logic_vector(to_unsigned( 20 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 112 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=818 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 82, 8)),
                    1 => std_logic_vector(to_unsigned( 29 , 8)),
                    2 => std_logic_vector(to_unsigned( 61 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 65 , 8)),
                    5 => std_logic_vector(to_unsigned( 14 , 8)),
                    6 => std_logic_vector(to_unsigned( 120 , 8)),
                    7 => std_logic_vector(to_unsigned( 105 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=819 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),
                    1 => std_logic_vector(to_unsigned( 84 , 8)),
                    2 => std_logic_vector(to_unsigned( 105 , 8)),
                    3 => std_logic_vector(to_unsigned( 101 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 109 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=820 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),
                    1 => std_logic_vector(to_unsigned( 84 , 8)),
                    2 => std_logic_vector(to_unsigned( 105 , 8)),
                    3 => std_logic_vector(to_unsigned( 101 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 109 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=821 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 115 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 68 , 8)),
                    4 => std_logic_vector(to_unsigned( 92 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 74 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=822 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 75 , 8)),
                    3 => std_logic_vector(to_unsigned( 110 , 8)),
                    4 => std_logic_vector(to_unsigned( 80 , 8)),
                    5 => std_logic_vector(to_unsigned( 7 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 99 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=823 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 75 , 8)),
                    3 => std_logic_vector(to_unsigned( 110 , 8)),
                    4 => std_logic_vector(to_unsigned( 80 , 8)),
                    5 => std_logic_vector(to_unsigned( 7 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 99 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=824 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 77, 8)),
                    1 => std_logic_vector(to_unsigned( 3 , 8)),
                    2 => std_logic_vector(to_unsigned( 82 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 60 , 8)),
                    5 => std_logic_vector(to_unsigned( 48 , 8)),
                    6 => std_logic_vector(to_unsigned( 93 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=825 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 56 , 8)),
                    3 => std_logic_vector(to_unsigned( 76 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 109 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=826 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 56 , 8)),
                    3 => std_logic_vector(to_unsigned( 76 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 109 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=827 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 26 , 8)),
                    2 => std_logic_vector(to_unsigned( 113 , 8)),
                    3 => std_logic_vector(to_unsigned( 118 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 58 , 8)),
                    7 => std_logic_vector(to_unsigned( 40 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=828 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),
                    1 => std_logic_vector(to_unsigned( 108 , 8)),
                    2 => std_logic_vector(to_unsigned( 11 , 8)),
                    3 => std_logic_vector(to_unsigned( 79 , 8)),
                    4 => std_logic_vector(to_unsigned( 57 , 8)),
                    5 => std_logic_vector(to_unsigned( 73 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 87 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=829 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),
                    1 => std_logic_vector(to_unsigned( 108 , 8)),
                    2 => std_logic_vector(to_unsigned( 11 , 8)),
                    3 => std_logic_vector(to_unsigned( 79 , 8)),
                    4 => std_logic_vector(to_unsigned( 57 , 8)),
                    5 => std_logic_vector(to_unsigned( 73 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 87 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=830 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 52 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 12 , 8)),
                    6 => std_logic_vector(to_unsigned( 63 , 8)),
                    7 => std_logic_vector(to_unsigned( 23 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=831 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 101 , 8)),
                    3 => std_logic_vector(to_unsigned( 65 , 8)),
                    4 => std_logic_vector(to_unsigned( 69 , 8)),
                    5 => std_logic_vector(to_unsigned( 105 , 8)),
                    6 => std_logic_vector(to_unsigned( 22 , 8)),
                    7 => std_logic_vector(to_unsigned( 17 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=832 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 101 , 8)),
                    3 => std_logic_vector(to_unsigned( 65 , 8)),
                    4 => std_logic_vector(to_unsigned( 69 , 8)),
                    5 => std_logic_vector(to_unsigned( 105 , 8)),
                    6 => std_logic_vector(to_unsigned( 22 , 8)),
                    7 => std_logic_vector(to_unsigned( 17 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=833 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),
                    1 => std_logic_vector(to_unsigned( 0 , 8)),
                    2 => std_logic_vector(to_unsigned( 87 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 116 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 91 , 8)),
                    7 => std_logic_vector(to_unsigned( 81 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=834 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 47 , 8)),
                    2 => std_logic_vector(to_unsigned( 38 , 8)),
                    3 => std_logic_vector(to_unsigned( 123 , 8)),
                    4 => std_logic_vector(to_unsigned( 23 , 8)),
                    5 => std_logic_vector(to_unsigned( 1 , 8)),
                    6 => std_logic_vector(to_unsigned( 68 , 8)),
                    7 => std_logic_vector(to_unsigned( 51 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=835 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 47 , 8)),
                    2 => std_logic_vector(to_unsigned( 38 , 8)),
                    3 => std_logic_vector(to_unsigned( 123 , 8)),
                    4 => std_logic_vector(to_unsigned( 23 , 8)),
                    5 => std_logic_vector(to_unsigned( 1 , 8)),
                    6 => std_logic_vector(to_unsigned( 68 , 8)),
                    7 => std_logic_vector(to_unsigned( 51 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=836 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),
                    1 => std_logic_vector(to_unsigned( 2 , 8)),
                    2 => std_logic_vector(to_unsigned( 51 , 8)),
                    3 => std_logic_vector(to_unsigned( 35 , 8)),
                    4 => std_logic_vector(to_unsigned( 59 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 78 , 8)),
                    7 => std_logic_vector(to_unsigned( 39 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=837 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 111 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 64 , 8)),
                    5 => std_logic_vector(to_unsigned( 36 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=838 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 111 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 64 , 8)),
                    5 => std_logic_vector(to_unsigned( 36 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=839 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),
                    1 => std_logic_vector(to_unsigned( 95 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 43 , 8)),
                    4 => std_logic_vector(to_unsigned( 83 , 8)),
                    5 => std_logic_vector(to_unsigned( 112 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 36 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=840 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 90 , 8)),
                    3 => std_logic_vector(to_unsigned( 39 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 29 , 8)),
                    6 => std_logic_vector(to_unsigned( 3 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=841 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 90 , 8)),
                    3 => std_logic_vector(to_unsigned( 39 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 29 , 8)),
                    6 => std_logic_vector(to_unsigned( 3 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=842 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 45 , 8)),
                    4 => std_logic_vector(to_unsigned( 106 , 8)),
                    5 => std_logic_vector(to_unsigned( 34 , 8)),
                    6 => std_logic_vector(to_unsigned( 51 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=843 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 63, 8)),
                    1 => std_logic_vector(to_unsigned( 92 , 8)),
                    2 => std_logic_vector(to_unsigned( 104 , 8)),
                    3 => std_logic_vector(to_unsigned( 8 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 12 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=844 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 63, 8)),
                    1 => std_logic_vector(to_unsigned( 92 , 8)),
                    2 => std_logic_vector(to_unsigned( 104 , 8)),
                    3 => std_logic_vector(to_unsigned( 8 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 12 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=845 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 33, 8)),
                    1 => std_logic_vector(to_unsigned( 10 , 8)),
                    2 => std_logic_vector(to_unsigned( 47 , 8)),
                    3 => std_logic_vector(to_unsigned( 28 , 8)),
                    4 => std_logic_vector(to_unsigned( 14 , 8)),
                    5 => std_logic_vector(to_unsigned( 82 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 76 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=846 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),
                    1 => std_logic_vector(to_unsigned( 103 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 63 , 8)),
                    4 => std_logic_vector(to_unsigned( 114 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 110 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=847 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),
                    1 => std_logic_vector(to_unsigned( 103 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 63 , 8)),
                    4 => std_logic_vector(to_unsigned( 114 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 110 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=848 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),
                    1 => std_logic_vector(to_unsigned( 94 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 23 , 8)),
                    4 => std_logic_vector(to_unsigned( 98 , 8)),
                    5 => std_logic_vector(to_unsigned( 120 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 103 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=849 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),
                    1 => std_logic_vector(to_unsigned( 24 , 8)),
                    2 => std_logic_vector(to_unsigned( 81 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 96 , 8)),
                    5 => std_logic_vector(to_unsigned( 5 , 8)),
                    6 => std_logic_vector(to_unsigned( 59 , 8)),
                    7 => std_logic_vector(to_unsigned( 69 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=850 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),
                    1 => std_logic_vector(to_unsigned( 24 , 8)),
                    2 => std_logic_vector(to_unsigned( 81 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 96 , 8)),
                    5 => std_logic_vector(to_unsigned( 5 , 8)),
                    6 => std_logic_vector(to_unsigned( 59 , 8)),
                    7 => std_logic_vector(to_unsigned( 69 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=851 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 109, 8)),
                    1 => std_logic_vector(to_unsigned( 123 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 65 , 8)),
                    4 => std_logic_vector(to_unsigned( 49 , 8)),
                    5 => std_logic_vector(to_unsigned( 72 , 8)),
                    6 => std_logic_vector(to_unsigned( 32 , 8)),
                    7 => std_logic_vector(to_unsigned( 39 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=852 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 80, 8)),
                    1 => std_logic_vector(to_unsigned( 123 , 8)),
                    2 => std_logic_vector(to_unsigned( 106 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 24 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 52 , 8)),
                    7 => std_logic_vector(to_unsigned( 110 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=853 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 80, 8)),
                    1 => std_logic_vector(to_unsigned( 123 , 8)),
                    2 => std_logic_vector(to_unsigned( 106 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 24 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 52 , 8)),
                    7 => std_logic_vector(to_unsigned( 110 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=854 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 47, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 9 , 8)),
                    3 => std_logic_vector(to_unsigned( 84 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 56 , 8)),
                    6 => std_logic_vector(to_unsigned( 74 , 8)),
                    7 => std_logic_vector(to_unsigned( 98 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=855 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 96, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 30 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 116 , 8)),
                    5 => std_logic_vector(to_unsigned( 48 , 8)),
                    6 => std_logic_vector(to_unsigned( 8 , 8)),
                    7 => std_logic_vector(to_unsigned( 71 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=856 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 96, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 30 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 116 , 8)),
                    5 => std_logic_vector(to_unsigned( 48 , 8)),
                    6 => std_logic_vector(to_unsigned( 8 , 8)),
                    7 => std_logic_vector(to_unsigned( 71 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=857 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 99, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 39 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 61 , 8)),
                    6 => std_logic_vector(to_unsigned( 2 , 8)),
                    7 => std_logic_vector(to_unsigned( 68 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=858 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),
                    1 => std_logic_vector(to_unsigned( 39 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 8 , 8)),
                    4 => std_logic_vector(to_unsigned( 59 , 8)),
                    5 => std_logic_vector(to_unsigned( 45 , 8)),
                    6 => std_logic_vector(to_unsigned( 31 , 8)),
                    7 => std_logic_vector(to_unsigned( 97 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=859 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),
                    1 => std_logic_vector(to_unsigned( 39 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 8 , 8)),
                    4 => std_logic_vector(to_unsigned( 59 , 8)),
                    5 => std_logic_vector(to_unsigned( 45 , 8)),
                    6 => std_logic_vector(to_unsigned( 31 , 8)),
                    7 => std_logic_vector(to_unsigned( 97 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=860 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),
                    1 => std_logic_vector(to_unsigned( 56 , 8)),
                    2 => std_logic_vector(to_unsigned( 28 , 8)),
                    3 => std_logic_vector(to_unsigned( 49 , 8)),
                    4 => std_logic_vector(to_unsigned( 3 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 105 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=861 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 33, 8)),
                    1 => std_logic_vector(to_unsigned( 65 , 8)),
                    2 => std_logic_vector(to_unsigned( 90 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 27 , 8)),
                    5 => std_logic_vector(to_unsigned( 10 , 8)),
                    6 => std_logic_vector(to_unsigned( 115 , 8)),
                    7 => std_logic_vector(to_unsigned( 48 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=862 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 33, 8)),
                    1 => std_logic_vector(to_unsigned( 65 , 8)),
                    2 => std_logic_vector(to_unsigned( 90 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 27 , 8)),
                    5 => std_logic_vector(to_unsigned( 10 , 8)),
                    6 => std_logic_vector(to_unsigned( 115 , 8)),
                    7 => std_logic_vector(to_unsigned( 48 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=863 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 87 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 47 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 39 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=864 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 67 , 8)),
                    2 => std_logic_vector(to_unsigned( 60 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 42 , 8)),
                    5 => std_logic_vector(to_unsigned( 37 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=865 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 67 , 8)),
                    2 => std_logic_vector(to_unsigned( 60 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 42 , 8)),
                    5 => std_logic_vector(to_unsigned( 37 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=866 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),
                    1 => std_logic_vector(to_unsigned( 12 , 8)),
                    2 => std_logic_vector(to_unsigned( 79 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 57 , 8)),
                    5 => std_logic_vector(to_unsigned( 68 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 45 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=867 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 9 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 117 , 8)),
                    6 => std_logic_vector(to_unsigned( 97 , 8)),
                    7 => std_logic_vector(to_unsigned( 1 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=868 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 9 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 117 , 8)),
                    6 => std_logic_vector(to_unsigned( 97 , 8)),
                    7 => std_logic_vector(to_unsigned( 1 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=869 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 70, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 38 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 118 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 15 , 8)),
                    7 => std_logic_vector(to_unsigned( 10 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=870 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),
                    1 => std_logic_vector(to_unsigned( 61 , 8)),
                    2 => std_logic_vector(to_unsigned( 100 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 123 , 8)),
                    6 => std_logic_vector(to_unsigned( 32 , 8)),
                    7 => std_logic_vector(to_unsigned( 8 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=871 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),
                    1 => std_logic_vector(to_unsigned( 61 , 8)),
                    2 => std_logic_vector(to_unsigned( 100 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 123 , 8)),
                    6 => std_logic_vector(to_unsigned( 32 , 8)),
                    7 => std_logic_vector(to_unsigned( 8 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=872 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 40, 8)),
                    1 => std_logic_vector(to_unsigned( 71 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 59 , 8)),
                    4 => std_logic_vector(to_unsigned( 24 , 8)),
                    5 => std_logic_vector(to_unsigned( 100 , 8)),
                    6 => std_logic_vector(to_unsigned( 28 , 8)),
                    7 => std_logic_vector(to_unsigned( 117 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=873 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 91, 8)),
                    1 => std_logic_vector(to_unsigned( 17 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 86 , 8)),
                    4 => std_logic_vector(to_unsigned( 121 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 66 , 8)),
                    7 => std_logic_vector(to_unsigned( 116 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=874 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 91, 8)),
                    1 => std_logic_vector(to_unsigned( 17 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 86 , 8)),
                    4 => std_logic_vector(to_unsigned( 121 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 66 , 8)),
                    7 => std_logic_vector(to_unsigned( 116 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=875 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 20, 8)),
                    1 => std_logic_vector(to_unsigned( 119 , 8)),
                    2 => std_logic_vector(to_unsigned( 105 , 8)),
                    3 => std_logic_vector(to_unsigned( 5 , 8)),
                    4 => std_logic_vector(to_unsigned( 60 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 82 , 8)),
                    7 => std_logic_vector(to_unsigned( 69 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=876 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),
                    1 => std_logic_vector(to_unsigned( 50 , 8)),
                    2 => std_logic_vector(to_unsigned( 111 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 122 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 85 , 8)),
                    7 => std_logic_vector(to_unsigned( 28 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=877 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),
                    1 => std_logic_vector(to_unsigned( 50 , 8)),
                    2 => std_logic_vector(to_unsigned( 111 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 122 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 85 , 8)),
                    7 => std_logic_vector(to_unsigned( 28 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=878 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 67, 8)),
                    1 => std_logic_vector(to_unsigned( 72 , 8)),
                    2 => std_logic_vector(to_unsigned( 85 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 20 , 8)),
                    5 => std_logic_vector(to_unsigned( 62 , 8)),
                    6 => std_logic_vector(to_unsigned( 15 , 8)),
                    7 => std_logic_vector(to_unsigned( 98 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=879 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 40 , 8)),
                    2 => std_logic_vector(to_unsigned( 45 , 8)),
                    3 => std_logic_vector(to_unsigned( 7 , 8)),
                    4 => std_logic_vector(to_unsigned( 123 , 8)),
                    5 => std_logic_vector(to_unsigned( 90 , 8)),
                    6 => std_logic_vector(to_unsigned( 70 , 8)),
                    7 => std_logic_vector(to_unsigned( 78 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=880 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 40 , 8)),
                    2 => std_logic_vector(to_unsigned( 45 , 8)),
                    3 => std_logic_vector(to_unsigned( 7 , 8)),
                    4 => std_logic_vector(to_unsigned( 123 , 8)),
                    5 => std_logic_vector(to_unsigned( 90 , 8)),
                    6 => std_logic_vector(to_unsigned( 70 , 8)),
                    7 => std_logic_vector(to_unsigned( 78 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=881 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),
                    1 => std_logic_vector(to_unsigned( 33 , 8)),
                    2 => std_logic_vector(to_unsigned( 86 , 8)),
                    3 => std_logic_vector(to_unsigned( 124 , 8)),
                    4 => std_logic_vector(to_unsigned( 56 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 65 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=882 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),
                    1 => std_logic_vector(to_unsigned( 59 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 11 , 8)),
                    5 => std_logic_vector(to_unsigned( 75 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 111 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=883 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),
                    1 => std_logic_vector(to_unsigned( 59 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 11 , 8)),
                    5 => std_logic_vector(to_unsigned( 75 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 111 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=884 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 34 , 8)),
                    3 => std_logic_vector(to_unsigned( 66 , 8)),
                    4 => std_logic_vector(to_unsigned( 116 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=885 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 98 , 8)),
                    3 => std_logic_vector(to_unsigned( 28 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 55 , 8)),
                    6 => std_logic_vector(to_unsigned( 33 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=886 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 98 , 8)),
                    3 => std_logic_vector(to_unsigned( 28 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 55 , 8)),
                    6 => std_logic_vector(to_unsigned( 33 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=887 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 113, 8)),
                    1 => std_logic_vector(to_unsigned( 75 , 8)),
                    2 => std_logic_vector(to_unsigned( 32 , 8)),
                    3 => std_logic_vector(to_unsigned( 12 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 50 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=888 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 20, 8)),
                    1 => std_logic_vector(to_unsigned( 112 , 8)),
                    2 => std_logic_vector(to_unsigned( 63 , 8)),
                    3 => std_logic_vector(to_unsigned( 25 , 8)),
                    4 => std_logic_vector(to_unsigned( 69 , 8)),
                    5 => std_logic_vector(to_unsigned( 92 , 8)),
                    6 => std_logic_vector(to_unsigned( 106 , 8)),
                    7 => std_logic_vector(to_unsigned( 116 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=889 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 20, 8)),
                    1 => std_logic_vector(to_unsigned( 112 , 8)),
                    2 => std_logic_vector(to_unsigned( 63 , 8)),
                    3 => std_logic_vector(to_unsigned( 25 , 8)),
                    4 => std_logic_vector(to_unsigned( 69 , 8)),
                    5 => std_logic_vector(to_unsigned( 92 , 8)),
                    6 => std_logic_vector(to_unsigned( 106 , 8)),
                    7 => std_logic_vector(to_unsigned( 116 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=890 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 69 , 8)),
                    4 => std_logic_vector(to_unsigned( 63 , 8)),
                    5 => std_logic_vector(to_unsigned( 47 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=891 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),
                    1 => std_logic_vector(to_unsigned( 63 , 8)),
                    2 => std_logic_vector(to_unsigned( 117 , 8)),
                    3 => std_logic_vector(to_unsigned( 28 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 105 , 8)),
                    6 => std_logic_vector(to_unsigned( 7 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=892 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),
                    1 => std_logic_vector(to_unsigned( 63 , 8)),
                    2 => std_logic_vector(to_unsigned( 117 , 8)),
                    3 => std_logic_vector(to_unsigned( 28 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 105 , 8)),
                    6 => std_logic_vector(to_unsigned( 7 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=893 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 111 , 8)),
                    3 => std_logic_vector(to_unsigned( 86 , 8)),
                    4 => std_logic_vector(to_unsigned( 39 , 8)),
                    5 => std_logic_vector(to_unsigned( 6 , 8)),
                    6 => std_logic_vector(to_unsigned( 35 , 8)),
                    7 => std_logic_vector(to_unsigned( 18 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=894 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 95 , 8)),
                    4 => std_logic_vector(to_unsigned( 9 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 39 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=895 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 95 , 8)),
                    4 => std_logic_vector(to_unsigned( 9 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 39 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=896 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 23 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 124 , 8)),
                    6 => std_logic_vector(to_unsigned( 69 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=897 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 2 , 8)),
                    2 => std_logic_vector(to_unsigned( 49 , 8)),
                    3 => std_logic_vector(to_unsigned( 115 , 8)),
                    4 => std_logic_vector(to_unsigned( 82 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 35 , 8)),
                    7 => std_logic_vector(to_unsigned( 64 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=898 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 2 , 8)),
                    2 => std_logic_vector(to_unsigned( 49 , 8)),
                    3 => std_logic_vector(to_unsigned( 115 , 8)),
                    4 => std_logic_vector(to_unsigned( 82 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 35 , 8)),
                    7 => std_logic_vector(to_unsigned( 64 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=899 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 118, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 83 , 8)),
                    3 => std_logic_vector(to_unsigned( 71 , 8)),
                    4 => std_logic_vector(to_unsigned( 40 , 8)),
                    5 => std_logic_vector(to_unsigned( 56 , 8)),
                    6 => std_logic_vector(to_unsigned( 67 , 8)),
                    7 => std_logic_vector(to_unsigned( 107 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=900 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 100 , 8)),
                    2 => std_logic_vector(to_unsigned( 109 , 8)),
                    3 => std_logic_vector(to_unsigned( 56 , 8)),
                    4 => std_logic_vector(to_unsigned( 40 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 78 , 8)),
                    7 => std_logic_vector(to_unsigned( 18 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=901 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 100 , 8)),
                    2 => std_logic_vector(to_unsigned( 109 , 8)),
                    3 => std_logic_vector(to_unsigned( 56 , 8)),
                    4 => std_logic_vector(to_unsigned( 40 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 78 , 8)),
                    7 => std_logic_vector(to_unsigned( 18 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=902 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 94, 8)),
                    1 => std_logic_vector(to_unsigned( 21 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 26 , 8)),
                    4 => std_logic_vector(to_unsigned( 51 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 82 , 8)),
                    7 => std_logic_vector(to_unsigned( 55 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=903 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 38 , 8)),
                    2 => std_logic_vector(to_unsigned( 42 , 8)),
                    3 => std_logic_vector(to_unsigned( 110 , 8)),
                    4 => std_logic_vector(to_unsigned( 97 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 58 , 8)),
                    7 => std_logic_vector(to_unsigned( 22 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=904 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 38 , 8)),
                    2 => std_logic_vector(to_unsigned( 42 , 8)),
                    3 => std_logic_vector(to_unsigned( 110 , 8)),
                    4 => std_logic_vector(to_unsigned( 97 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 58 , 8)),
                    7 => std_logic_vector(to_unsigned( 22 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=905 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 115, 8)),
                    1 => std_logic_vector(to_unsigned( 59 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 99 , 8)),
                    4 => std_logic_vector(to_unsigned( 2 , 8)),
                    5 => std_logic_vector(to_unsigned( 87 , 8)),
                    6 => std_logic_vector(to_unsigned( 14 , 8)),
                    7 => std_logic_vector(to_unsigned( 107 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=906 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 25, 8)),
                    1 => std_logic_vector(to_unsigned( 65 , 8)),
                    2 => std_logic_vector(to_unsigned( 86 , 8)),
                    3 => std_logic_vector(to_unsigned( 112 , 8)),
                    4 => std_logic_vector(to_unsigned( 97 , 8)),
                    5 => std_logic_vector(to_unsigned( 124 , 8)),
                    6 => std_logic_vector(to_unsigned( 20 , 8)),
                    7 => std_logic_vector(to_unsigned( 42 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=907 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 25, 8)),
                    1 => std_logic_vector(to_unsigned( 65 , 8)),
                    2 => std_logic_vector(to_unsigned( 86 , 8)),
                    3 => std_logic_vector(to_unsigned( 112 , 8)),
                    4 => std_logic_vector(to_unsigned( 97 , 8)),
                    5 => std_logic_vector(to_unsigned( 124 , 8)),
                    6 => std_logic_vector(to_unsigned( 20 , 8)),
                    7 => std_logic_vector(to_unsigned( 42 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=908 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 88, 8)),
                    1 => std_logic_vector(to_unsigned( 33 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 44 , 8)),
                    4 => std_logic_vector(to_unsigned( 51 , 8)),
                    5 => std_logic_vector(to_unsigned( 20 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 108 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=909 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 53 , 8)),
                    3 => std_logic_vector(to_unsigned( 49 , 8)),
                    4 => std_logic_vector(to_unsigned( 23 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 1 , 8)),
                    7 => std_logic_vector(to_unsigned( 77 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=910 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 53 , 8)),
                    3 => std_logic_vector(to_unsigned( 49 , 8)),
                    4 => std_logic_vector(to_unsigned( 23 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 1 , 8)),
                    7 => std_logic_vector(to_unsigned( 77 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=911 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),
                    1 => std_logic_vector(to_unsigned( 120 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 105 , 8)),
                    5 => std_logic_vector(to_unsigned( 61 , 8)),
                    6 => std_logic_vector(to_unsigned( 57 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=912 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 118, 8)),
                    1 => std_logic_vector(to_unsigned( 39 , 8)),
                    2 => std_logic_vector(to_unsigned( 34 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 67 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 30 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=913 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 118, 8)),
                    1 => std_logic_vector(to_unsigned( 39 , 8)),
                    2 => std_logic_vector(to_unsigned( 34 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 67 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 30 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=914 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),
                    1 => std_logic_vector(to_unsigned( 99 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 44 , 8)),
                    4 => std_logic_vector(to_unsigned( 10 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 32 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=915 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 98 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 72 , 8)),
                    5 => std_logic_vector(to_unsigned( 76 , 8)),
                    6 => std_logic_vector(to_unsigned( 44 , 8)),
                    7 => std_logic_vector(to_unsigned( 56 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=916 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 98 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 72 , 8)),
                    5 => std_logic_vector(to_unsigned( 76 , 8)),
                    6 => std_logic_vector(to_unsigned( 44 , 8)),
                    7 => std_logic_vector(to_unsigned( 56 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=917 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 33, 8)),
                    1 => std_logic_vector(to_unsigned( 121 , 8)),
                    2 => std_logic_vector(to_unsigned( 75 , 8)),
                    3 => std_logic_vector(to_unsigned( 86 , 8)),
                    4 => std_logic_vector(to_unsigned( 40 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 114 , 8)),
                    7 => std_logic_vector(to_unsigned( 60 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=918 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 42 , 8)),
                    3 => std_logic_vector(to_unsigned( 11 , 8)),
                    4 => std_logic_vector(to_unsigned( 97 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 93 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=919 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 42 , 8)),
                    3 => std_logic_vector(to_unsigned( 11 , 8)),
                    4 => std_logic_vector(to_unsigned( 97 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 93 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=920 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),
                    1 => std_logic_vector(to_unsigned( 46 , 8)),
                    2 => std_logic_vector(to_unsigned( 36 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 83 , 8)),
                    5 => std_logic_vector(to_unsigned( 112 , 8)),
                    6 => std_logic_vector(to_unsigned( 104 , 8)),
                    7 => std_logic_vector(to_unsigned( 118 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=921 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),
                    1 => std_logic_vector(to_unsigned( 103 , 8)),
                    2 => std_logic_vector(to_unsigned( 60 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 6 , 8)),
                    6 => std_logic_vector(to_unsigned( 69 , 8)),
                    7 => std_logic_vector(to_unsigned( 11 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=922 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),
                    1 => std_logic_vector(to_unsigned( 103 , 8)),
                    2 => std_logic_vector(to_unsigned( 60 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 6 , 8)),
                    6 => std_logic_vector(to_unsigned( 69 , 8)),
                    7 => std_logic_vector(to_unsigned( 11 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=923 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),
                    1 => std_logic_vector(to_unsigned( 107 , 8)),
                    2 => std_logic_vector(to_unsigned( 122 , 8)),
                    3 => std_logic_vector(to_unsigned( 39 , 8)),
                    4 => std_logic_vector(to_unsigned( 93 , 8)),
                    5 => std_logic_vector(to_unsigned( 77 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=924 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),
                    1 => std_logic_vector(to_unsigned( 86 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 98 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 82 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 55 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=925 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),
                    1 => std_logic_vector(to_unsigned( 86 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 98 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 82 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 55 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=926 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 114 , 8)),
                    3 => std_logic_vector(to_unsigned( 102 , 8)),
                    4 => std_logic_vector(to_unsigned( 31 , 8)),
                    5 => std_logic_vector(to_unsigned( 119 , 8)),
                    6 => std_logic_vector(to_unsigned( 14 , 8)),
                    7 => std_logic_vector(to_unsigned( 21 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=927 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 110, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 1 , 8)),
                    3 => std_logic_vector(to_unsigned( 104 , 8)),
                    4 => std_logic_vector(to_unsigned( 31 , 8)),
                    5 => std_logic_vector(to_unsigned( 52 , 8)),
                    6 => std_logic_vector(to_unsigned( 16 , 8)),
                    7 => std_logic_vector(to_unsigned( 68 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=928 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 110, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 1 , 8)),
                    3 => std_logic_vector(to_unsigned( 104 , 8)),
                    4 => std_logic_vector(to_unsigned( 31 , 8)),
                    5 => std_logic_vector(to_unsigned( 52 , 8)),
                    6 => std_logic_vector(to_unsigned( 16 , 8)),
                    7 => std_logic_vector(to_unsigned( 68 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=929 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 83, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 68 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 0 , 8)),
                    6 => std_logic_vector(to_unsigned( 42 , 8)),
                    7 => std_logic_vector(to_unsigned( 19 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=930 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 12, 8)),
                    1 => std_logic_vector(to_unsigned( 81 , 8)),
                    2 => std_logic_vector(to_unsigned( 56 , 8)),
                    3 => std_logic_vector(to_unsigned( 69 , 8)),
                    4 => std_logic_vector(to_unsigned( 120 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 110 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=931 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 12, 8)),
                    1 => std_logic_vector(to_unsigned( 81 , 8)),
                    2 => std_logic_vector(to_unsigned( 56 , 8)),
                    3 => std_logic_vector(to_unsigned( 69 , 8)),
                    4 => std_logic_vector(to_unsigned( 120 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 110 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=932 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),
                    1 => std_logic_vector(to_unsigned( 77 , 8)),
                    2 => std_logic_vector(to_unsigned( 22 , 8)),
                    3 => std_logic_vector(to_unsigned( 96 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 112 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=933 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 120 , 8)),
                    3 => std_logic_vector(to_unsigned( 66 , 8)),
                    4 => std_logic_vector(to_unsigned( 98 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 57 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=934 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 120 , 8)),
                    3 => std_logic_vector(to_unsigned( 66 , 8)),
                    4 => std_logic_vector(to_unsigned( 98 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 57 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=935 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),
                    1 => std_logic_vector(to_unsigned( 108 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 103 , 8)),
                    4 => std_logic_vector(to_unsigned( 80 , 8)),
                    5 => std_logic_vector(to_unsigned( 25 , 8)),
                    6 => std_logic_vector(to_unsigned( 73 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=936 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),
                    1 => std_logic_vector(to_unsigned( 35 , 8)),
                    2 => std_logic_vector(to_unsigned( 78 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 101 , 8)),
                    5 => std_logic_vector(to_unsigned( 11 , 8)),
                    6 => std_logic_vector(to_unsigned( 41 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=937 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),
                    1 => std_logic_vector(to_unsigned( 35 , 8)),
                    2 => std_logic_vector(to_unsigned( 78 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 101 , 8)),
                    5 => std_logic_vector(to_unsigned( 11 , 8)),
                    6 => std_logic_vector(to_unsigned( 41 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=938 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 97, 8)),
                    1 => std_logic_vector(to_unsigned( 71 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 30 , 8)),
                    6 => std_logic_vector(to_unsigned( 21 , 8)),
                    7 => std_logic_vector(to_unsigned( 14 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=939 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 108 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 39 , 8)),
                    6 => std_logic_vector(to_unsigned( 123 , 8)),
                    7 => std_logic_vector(to_unsigned( 58 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=940 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 108 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 39 , 8)),
                    6 => std_logic_vector(to_unsigned( 123 , 8)),
                    7 => std_logic_vector(to_unsigned( 58 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=941 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 109, 8)),
                    1 => std_logic_vector(to_unsigned( 51 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 96 , 8)),
                    4 => std_logic_vector(to_unsigned( 40 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 14 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=942 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 92 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 45 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 124 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=943 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 92 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 45 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 124 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=944 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 65 , 8)),
                    2 => std_logic_vector(to_unsigned( 37 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 31 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 114 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=945 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),
                    1 => std_logic_vector(to_unsigned( 25 , 8)),
                    2 => std_logic_vector(to_unsigned( 98 , 8)),
                    3 => std_logic_vector(to_unsigned( 7 , 8)),
                    4 => std_logic_vector(to_unsigned( 94 , 8)),
                    5 => std_logic_vector(to_unsigned( 88 , 8)),
                    6 => std_logic_vector(to_unsigned( 82 , 8)),
                    7 => std_logic_vector(to_unsigned( 104 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=946 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),
                    1 => std_logic_vector(to_unsigned( 25 , 8)),
                    2 => std_logic_vector(to_unsigned( 98 , 8)),
                    3 => std_logic_vector(to_unsigned( 7 , 8)),
                    4 => std_logic_vector(to_unsigned( 94 , 8)),
                    5 => std_logic_vector(to_unsigned( 88 , 8)),
                    6 => std_logic_vector(to_unsigned( 82 , 8)),
                    7 => std_logic_vector(to_unsigned( 104 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=947 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 108 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 24 , 8)),
                    6 => std_logic_vector(to_unsigned( 67 , 8)),
                    7 => std_logic_vector(to_unsigned( 94 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=948 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 17, 8)),
                    1 => std_logic_vector(to_unsigned( 118 , 8)),
                    2 => std_logic_vector(to_unsigned( 104 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 40 , 8)),
                    5 => std_logic_vector(to_unsigned( 54 , 8)),
                    6 => std_logic_vector(to_unsigned( 48 , 8)),
                    7 => std_logic_vector(to_unsigned( 83 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=949 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 17, 8)),
                    1 => std_logic_vector(to_unsigned( 118 , 8)),
                    2 => std_logic_vector(to_unsigned( 104 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 40 , 8)),
                    5 => std_logic_vector(to_unsigned( 54 , 8)),
                    6 => std_logic_vector(to_unsigned( 48 , 8)),
                    7 => std_logic_vector(to_unsigned( 83 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=950 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 16, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 88 , 8)),
                    3 => std_logic_vector(to_unsigned( 119 , 8)),
                    4 => std_logic_vector(to_unsigned( 54 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 113 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=951 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 90 , 8)),
                    3 => std_logic_vector(to_unsigned( 82 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 121 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=952 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 90 , 8)),
                    3 => std_logic_vector(to_unsigned( 82 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 121 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=953 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 114 , 8)),
                    3 => std_logic_vector(to_unsigned( 103 , 8)),
                    4 => std_logic_vector(to_unsigned( 93 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 56 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=954 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 8, 8)),
                    1 => std_logic_vector(to_unsigned( 103 , 8)),
                    2 => std_logic_vector(to_unsigned( 80 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 4 , 8)),
                    5 => std_logic_vector(to_unsigned( 21 , 8)),
                    6 => std_logic_vector(to_unsigned( 65 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=955 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 8, 8)),
                    1 => std_logic_vector(to_unsigned( 103 , 8)),
                    2 => std_logic_vector(to_unsigned( 80 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 4 , 8)),
                    5 => std_logic_vector(to_unsigned( 21 , 8)),
                    6 => std_logic_vector(to_unsigned( 65 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=956 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 86 , 8)),
                    2 => std_logic_vector(to_unsigned( 68 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 24 , 8)),
                    5 => std_logic_vector(to_unsigned( 49 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=957 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 16, 8)),
                    1 => std_logic_vector(to_unsigned( 39 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 67 , 8)),
                    4 => std_logic_vector(to_unsigned( 75 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 85 , 8)),
                    7 => std_logic_vector(to_unsigned( 56 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=958 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 16, 8)),
                    1 => std_logic_vector(to_unsigned( 39 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 67 , 8)),
                    4 => std_logic_vector(to_unsigned( 75 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 85 , 8)),
                    7 => std_logic_vector(to_unsigned( 56 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=959 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 113, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 19 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 84 , 8)),
                    6 => std_logic_vector(to_unsigned( 92 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=960 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 90 , 8)),
                    2 => std_logic_vector(to_unsigned( 71 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 101 , 8)),
                    6 => std_logic_vector(to_unsigned( 65 , 8)),
                    7 => std_logic_vector(to_unsigned( 16 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=961 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 90 , 8)),
                    2 => std_logic_vector(to_unsigned( 71 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 101 , 8)),
                    6 => std_logic_vector(to_unsigned( 65 , 8)),
                    7 => std_logic_vector(to_unsigned( 16 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=962 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 12, 8)),
                    1 => std_logic_vector(to_unsigned( 99 , 8)),
                    2 => std_logic_vector(to_unsigned( 68 , 8)),
                    3 => std_logic_vector(to_unsigned( 84 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 7 , 8)),
                    6 => std_logic_vector(to_unsigned( 121 , 8)),
                    7 => std_logic_vector(to_unsigned( 53 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=963 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 37 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 82 , 8)),
                    5 => std_logic_vector(to_unsigned( 122 , 8)),
                    6 => std_logic_vector(to_unsigned( 52 , 8)),
                    7 => std_logic_vector(to_unsigned( 101 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=964 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 37 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 82 , 8)),
                    5 => std_logic_vector(to_unsigned( 122 , 8)),
                    6 => std_logic_vector(to_unsigned( 52 , 8)),
                    7 => std_logic_vector(to_unsigned( 101 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=965 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 21 , 8)),
                    2 => std_logic_vector(to_unsigned( 115 , 8)),
                    3 => std_logic_vector(to_unsigned( 88 , 8)),
                    4 => std_logic_vector(to_unsigned( 97 , 8)),
                    5 => std_logic_vector(to_unsigned( 43 , 8)),
                    6 => std_logic_vector(to_unsigned( 1 , 8)),
                    7 => std_logic_vector(to_unsigned( 74 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=966 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 120 , 8)),
                    2 => std_logic_vector(to_unsigned( 71 , 8)),
                    3 => std_logic_vector(to_unsigned( 67 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 35 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=967 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 120 , 8)),
                    2 => std_logic_vector(to_unsigned( 71 , 8)),
                    3 => std_logic_vector(to_unsigned( 67 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 35 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=968 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),
                    1 => std_logic_vector(to_unsigned( 44 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 21 , 8)),
                    4 => std_logic_vector(to_unsigned( 8 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 29 , 8)),
                    7 => std_logic_vector(to_unsigned( 83 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=969 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 105 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 17 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=970 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 105 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 17 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=971 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 66 , 8)),
                    2 => std_logic_vector(to_unsigned( 36 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 21 , 8)),
                    5 => std_logic_vector(to_unsigned( 27 , 8)),
                    6 => std_logic_vector(to_unsigned( 42 , 8)),
                    7 => std_logic_vector(to_unsigned( 112 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=972 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 38, 8)),
                    1 => std_logic_vector(to_unsigned( 63 , 8)),
                    2 => std_logic_vector(to_unsigned( 46 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 25 , 8)),
                    5 => std_logic_vector(to_unsigned( 54 , 8)),
                    6 => std_logic_vector(to_unsigned( 69 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=973 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 38, 8)),
                    1 => std_logic_vector(to_unsigned( 63 , 8)),
                    2 => std_logic_vector(to_unsigned( 46 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 25 , 8)),
                    5 => std_logic_vector(to_unsigned( 54 , 8)),
                    6 => std_logic_vector(to_unsigned( 69 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=974 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),
                    1 => std_logic_vector(to_unsigned( 18 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 117 , 8)),
                    4 => std_logic_vector(to_unsigned( 26 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=975 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),
                    1 => std_logic_vector(to_unsigned( 109 , 8)),
                    2 => std_logic_vector(to_unsigned( 43 , 8)),
                    3 => std_logic_vector(to_unsigned( 14 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 8 , 8)),
                    6 => std_logic_vector(to_unsigned( 74 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=976 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),
                    1 => std_logic_vector(to_unsigned( 109 , 8)),
                    2 => std_logic_vector(to_unsigned( 43 , 8)),
                    3 => std_logic_vector(to_unsigned( 14 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 8 , 8)),
                    6 => std_logic_vector(to_unsigned( 74 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=977 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 4, 8)),
                    1 => std_logic_vector(to_unsigned( 89 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 124 , 8)),
                    4 => std_logic_vector(to_unsigned( 33 , 8)),
                    5 => std_logic_vector(to_unsigned( 93 , 8)),
                    6 => std_logic_vector(to_unsigned( 102 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=978 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 94 , 8)),
                    2 => std_logic_vector(to_unsigned( 37 , 8)),
                    3 => std_logic_vector(to_unsigned( 28 , 8)),
                    4 => std_logic_vector(to_unsigned( 10 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 90 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=979 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 94 , 8)),
                    2 => std_logic_vector(to_unsigned( 37 , 8)),
                    3 => std_logic_vector(to_unsigned( 28 , 8)),
                    4 => std_logic_vector(to_unsigned( 10 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 90 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=980 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),
                    1 => std_logic_vector(to_unsigned( 91 , 8)),
                    2 => std_logic_vector(to_unsigned( 109 , 8)),
                    3 => std_logic_vector(to_unsigned( 45 , 8)),
                    4 => std_logic_vector(to_unsigned( 60 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 66 , 8)),
                    7 => std_logic_vector(to_unsigned( 4 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=981 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 84 , 8)),
                    2 => std_logic_vector(to_unsigned( 26 , 8)),
                    3 => std_logic_vector(to_unsigned( 65 , 8)),
                    4 => std_logic_vector(to_unsigned( 124 , 8)),
                    5 => std_logic_vector(to_unsigned( 109 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 19 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=982 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 84 , 8)),
                    2 => std_logic_vector(to_unsigned( 26 , 8)),
                    3 => std_logic_vector(to_unsigned( 65 , 8)),
                    4 => std_logic_vector(to_unsigned( 124 , 8)),
                    5 => std_logic_vector(to_unsigned( 109 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 19 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=983 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 102 , 8)),
                    3 => std_logic_vector(to_unsigned( 39 , 8)),
                    4 => std_logic_vector(to_unsigned( 86 , 8)),
                    5 => std_logic_vector(to_unsigned( 45 , 8)),
                    6 => std_logic_vector(to_unsigned( 121 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=984 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 39 , 8)),
                    3 => std_logic_vector(to_unsigned( 96 , 8)),
                    4 => std_logic_vector(to_unsigned( 70 , 8)),
                    5 => std_logic_vector(to_unsigned( 78 , 8)),
                    6 => std_logic_vector(to_unsigned( 104 , 8)),
                    7 => std_logic_vector(to_unsigned( 8 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=985 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 39 , 8)),
                    3 => std_logic_vector(to_unsigned( 96 , 8)),
                    4 => std_logic_vector(to_unsigned( 70 , 8)),
                    5 => std_logic_vector(to_unsigned( 78 , 8)),
                    6 => std_logic_vector(to_unsigned( 104 , 8)),
                    7 => std_logic_vector(to_unsigned( 8 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=986 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 2, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 74 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 10 , 8)),
                    7 => std_logic_vector(to_unsigned( 47 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=987 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 95 , 8)),
                    2 => std_logic_vector(to_unsigned( 46 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 24 , 8)),
                    5 => std_logic_vector(to_unsigned( 18 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=988 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 95 , 8)),
                    2 => std_logic_vector(to_unsigned( 46 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 24 , 8)),
                    5 => std_logic_vector(to_unsigned( 18 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=989 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 118, 8)),
                    1 => std_logic_vector(to_unsigned( 23 , 8)),
                    2 => std_logic_vector(to_unsigned( 73 , 8)),
                    3 => std_logic_vector(to_unsigned( 41 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 101 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 28 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=990 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 31 , 8)),
                    2 => std_logic_vector(to_unsigned( 106 , 8)),
                    3 => std_logic_vector(to_unsigned( 70 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 42 , 8)),
                    6 => std_logic_vector(to_unsigned( 51 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=991 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 31 , 8)),
                    2 => std_logic_vector(to_unsigned( 106 , 8)),
                    3 => std_logic_vector(to_unsigned( 70 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 42 , 8)),
                    6 => std_logic_vector(to_unsigned( 51 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=992 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 52 , 8)),
                    2 => std_logic_vector(to_unsigned( 48 , 8)),
                    3 => std_logic_vector(to_unsigned( 40 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 44 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=993 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 121 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 100 , 8)),
                    6 => std_logic_vector(to_unsigned( 1 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=994 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 121 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 100 , 8)),
                    6 => std_logic_vector(to_unsigned( 1 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=995 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 72, 8)),
                    1 => std_logic_vector(to_unsigned( 47 , 8)),
                    2 => std_logic_vector(to_unsigned( 38 , 8)),
                    3 => std_logic_vector(to_unsigned( 13 , 8)),
                    4 => std_logic_vector(to_unsigned( 65 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 4 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=996 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 99, 8)),
                    1 => std_logic_vector(to_unsigned( 32 , 8)),
                    2 => std_logic_vector(to_unsigned( 68 , 8)),
                    3 => std_logic_vector(to_unsigned( 20 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 109 , 8)),
                    6 => std_logic_vector(to_unsigned( 56 , 8)),
                    7 => std_logic_vector(to_unsigned( 25 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=997 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 99, 8)),
                    1 => std_logic_vector(to_unsigned( 32 , 8)),
                    2 => std_logic_vector(to_unsigned( 68 , 8)),
                    3 => std_logic_vector(to_unsigned( 20 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 109 , 8)),
                    6 => std_logic_vector(to_unsigned( 56 , 8)),
                    7 => std_logic_vector(to_unsigned( 25 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=998 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 123 , 8)),
                    2 => std_logic_vector(to_unsigned( 43 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 32 , 8)),
                    6 => std_logic_vector(to_unsigned( 27 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=999 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 33 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 86 , 8)),
                    5 => std_logic_vector(to_unsigned( 73 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 100 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1000 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 33 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 86 , 8)),
                    5 => std_logic_vector(to_unsigned( 73 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 100 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1001 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 21 , 8)),
                    4 => std_logic_vector(to_unsigned( 57 , 8)),
                    5 => std_logic_vector(to_unsigned( 33 , 8)),
                    6 => std_logic_vector(to_unsigned( 80 , 8)),
                    7 => std_logic_vector(to_unsigned( 94 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1002 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 15 , 8)),
                    3 => std_logic_vector(to_unsigned( 40 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 46 , 8)),
                    6 => std_logic_vector(to_unsigned( 121 , 8)),
                    7 => std_logic_vector(to_unsigned( 65 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1003 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 15 , 8)),
                    3 => std_logic_vector(to_unsigned( 40 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 46 , 8)),
                    6 => std_logic_vector(to_unsigned( 121 , 8)),
                    7 => std_logic_vector(to_unsigned( 65 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1004 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),
                    1 => std_logic_vector(to_unsigned( 60 , 8)),
                    2 => std_logic_vector(to_unsigned( 106 , 8)),
                    3 => std_logic_vector(to_unsigned( 99 , 8)),
                    4 => std_logic_vector(to_unsigned( 69 , 8)),
                    5 => std_logic_vector(to_unsigned( 6 , 8)),
                    6 => std_logic_vector(to_unsigned( 78 , 8)),
                    7 => std_logic_vector(to_unsigned( 30 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1005 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),
                    1 => std_logic_vector(to_unsigned( 10 , 8)),
                    2 => std_logic_vector(to_unsigned( 75 , 8)),
                    3 => std_logic_vector(to_unsigned( 91 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 60 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1006 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),
                    1 => std_logic_vector(to_unsigned( 10 , 8)),
                    2 => std_logic_vector(to_unsigned( 75 , 8)),
                    3 => std_logic_vector(to_unsigned( 91 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 60 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1007 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),
                    1 => std_logic_vector(to_unsigned( 6 , 8)),
                    2 => std_logic_vector(to_unsigned( 65 , 8)),
                    3 => std_logic_vector(to_unsigned( 82 , 8)),
                    4 => std_logic_vector(to_unsigned( 92 , 8)),
                    5 => std_logic_vector(to_unsigned( 30 , 8)),
                    6 => std_logic_vector(to_unsigned( 116 , 8)),
                    7 => std_logic_vector(to_unsigned( 51 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1008 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 110, 8)),
                    1 => std_logic_vector(to_unsigned( 30 , 8)),
                    2 => std_logic_vector(to_unsigned( 121 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 19 , 8)),
                    7 => std_logic_vector(to_unsigned( 61 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1009 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 110, 8)),
                    1 => std_logic_vector(to_unsigned( 30 , 8)),
                    2 => std_logic_vector(to_unsigned( 121 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 19 , 8)),
                    7 => std_logic_vector(to_unsigned( 61 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1010 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 40, 8)),
                    1 => std_logic_vector(to_unsigned( 19 , 8)),
                    2 => std_logic_vector(to_unsigned( 94 , 8)),
                    3 => std_logic_vector(to_unsigned( 10 , 8)),
                    4 => std_logic_vector(to_unsigned( 60 , 8)),
                    5 => std_logic_vector(to_unsigned( 120 , 8)),
                    6 => std_logic_vector(to_unsigned( 113 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1011 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 111 , 8)),
                    3 => std_logic_vector(to_unsigned( 60 , 8)),
                    4 => std_logic_vector(to_unsigned( 18 , 8)),
                    5 => std_logic_vector(to_unsigned( 23 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 33 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1012 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 111 , 8)),
                    3 => std_logic_vector(to_unsigned( 60 , 8)),
                    4 => std_logic_vector(to_unsigned( 18 , 8)),
                    5 => std_logic_vector(to_unsigned( 23 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 33 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1013 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 99, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 37 , 8)),
                    4 => std_logic_vector(to_unsigned( 33 , 8)),
                    5 => std_logic_vector(to_unsigned( 72 , 8)),
                    6 => std_logic_vector(to_unsigned( 94 , 8)),
                    7 => std_logic_vector(to_unsigned( 18 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1014 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),
                    1 => std_logic_vector(to_unsigned( 0 , 8)),
                    2 => std_logic_vector(to_unsigned( 117 , 8)),
                    3 => std_logic_vector(to_unsigned( 89 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 40 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1015 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),
                    1 => std_logic_vector(to_unsigned( 0 , 8)),
                    2 => std_logic_vector(to_unsigned( 117 , 8)),
                    3 => std_logic_vector(to_unsigned( 89 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 40 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1016 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 104 , 8)),
                    2 => std_logic_vector(to_unsigned( 1 , 8)),
                    3 => std_logic_vector(to_unsigned( 23 , 8)),
                    4 => std_logic_vector(to_unsigned( 85 , 8)),
                    5 => std_logic_vector(to_unsigned( 19 , 8)),
                    6 => std_logic_vector(to_unsigned( 28 , 8)),
                    7 => std_logic_vector(to_unsigned( 55 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1017 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 0 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 36 , 8)),
                    4 => std_logic_vector(to_unsigned( 17 , 8)),
                    5 => std_logic_vector(to_unsigned( 22 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 26 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1018 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 0 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 36 , 8)),
                    4 => std_logic_vector(to_unsigned( 17 , 8)),
                    5 => std_logic_vector(to_unsigned( 22 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 26 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1019 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 67, 8)),
                    1 => std_logic_vector(to_unsigned( 10 , 8)),
                    2 => std_logic_vector(to_unsigned( 102 , 8)),
                    3 => std_logic_vector(to_unsigned( 15 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 51 , 8)),
                    7 => std_logic_vector(to_unsigned( 4 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1020 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 54, 8)),
                    1 => std_logic_vector(to_unsigned( 46 , 8)),
                    2 => std_logic_vector(to_unsigned( 36 , 8)),
                    3 => std_logic_vector(to_unsigned( 116 , 8)),
                    4 => std_logic_vector(to_unsigned( 21 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 79 , 8)),
                    7 => std_logic_vector(to_unsigned( 4 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1021 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 54, 8)),
                    1 => std_logic_vector(to_unsigned( 46 , 8)),
                    2 => std_logic_vector(to_unsigned( 36 , 8)),
                    3 => std_logic_vector(to_unsigned( 116 , 8)),
                    4 => std_logic_vector(to_unsigned( 21 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 79 , 8)),
                    7 => std_logic_vector(to_unsigned( 4 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1022 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 53, 8)),
                    1 => std_logic_vector(to_unsigned( 60 , 8)),
                    2 => std_logic_vector(to_unsigned( 74 , 8)),
                    3 => std_logic_vector(to_unsigned( 92 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 21 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 3 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1023 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),
                    1 => std_logic_vector(to_unsigned( 0 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 68 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 43 , 8)),
                    6 => std_logic_vector(to_unsigned( 117 , 8)),
                    7 => std_logic_vector(to_unsigned( 87 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1024 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),
                    1 => std_logic_vector(to_unsigned( 0 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 68 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 43 , 8)),
                    6 => std_logic_vector(to_unsigned( 117 , 8)),
                    7 => std_logic_vector(to_unsigned( 87 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1025 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),
                    1 => std_logic_vector(to_unsigned( 98 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 113 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 55 , 8)),
                    6 => std_logic_vector(to_unsigned( 89 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1026 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 101 , 8)),
                    2 => std_logic_vector(to_unsigned( 70 , 8)),
                    3 => std_logic_vector(to_unsigned( 16 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 117 , 8)),
                    6 => std_logic_vector(to_unsigned( 24 , 8)),
                    7 => std_logic_vector(to_unsigned( 112 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1027 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 101 , 8)),
                    2 => std_logic_vector(to_unsigned( 70 , 8)),
                    3 => std_logic_vector(to_unsigned( 16 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 117 , 8)),
                    6 => std_logic_vector(to_unsigned( 24 , 8)),
                    7 => std_logic_vector(to_unsigned( 112 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1028 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),
                    1 => std_logic_vector(to_unsigned( 15 , 8)),
                    2 => std_logic_vector(to_unsigned( 52 , 8)),
                    3 => std_logic_vector(to_unsigned( 96 , 8)),
                    4 => std_logic_vector(to_unsigned( 8 , 8)),
                    5 => std_logic_vector(to_unsigned( 92 , 8)),
                    6 => std_logic_vector(to_unsigned( 122 , 8)),
                    7 => std_logic_vector(to_unsigned( 112 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1029 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 39 , 8)),
                    2 => std_logic_vector(to_unsigned( 87 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 103 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 50 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1030 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 39 , 8)),
                    2 => std_logic_vector(to_unsigned( 87 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 103 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 50 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1031 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 31 , 8)),
                    2 => std_logic_vector(to_unsigned( 61 , 8)),
                    3 => std_logic_vector(to_unsigned( 56 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 23 , 8)),
                    6 => std_logic_vector(to_unsigned( 51 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1032 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 110, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 85 , 8)),
                    3 => std_logic_vector(to_unsigned( 58 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 51 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 99 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1033 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 110, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 85 , 8)),
                    3 => std_logic_vector(to_unsigned( 58 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 51 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 99 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1034 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 108 , 8)),
                    2 => std_logic_vector(to_unsigned( 86 , 8)),
                    3 => std_logic_vector(to_unsigned( 15 , 8)),
                    4 => std_logic_vector(to_unsigned( 91 , 8)),
                    5 => std_logic_vector(to_unsigned( 63 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1035 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),
                    1 => std_logic_vector(to_unsigned( 89 , 8)),
                    2 => std_logic_vector(to_unsigned( 38 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 66 , 8)),
                    5 => std_logic_vector(to_unsigned( 71 , 8)),
                    6 => std_logic_vector(to_unsigned( 111 , 8)),
                    7 => std_logic_vector(to_unsigned( 10 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1036 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),
                    1 => std_logic_vector(to_unsigned( 89 , 8)),
                    2 => std_logic_vector(to_unsigned( 38 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 66 , 8)),
                    5 => std_logic_vector(to_unsigned( 71 , 8)),
                    6 => std_logic_vector(to_unsigned( 111 , 8)),
                    7 => std_logic_vector(to_unsigned( 10 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1037 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),
                    1 => std_logic_vector(to_unsigned( 80 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 92 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 5 , 8)),
                    6 => std_logic_vector(to_unsigned( 46 , 8)),
                    7 => std_logic_vector(to_unsigned( 108 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1038 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 111 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 115 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1039 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 111 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 115 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1040 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 70, 8)),
                    1 => std_logic_vector(to_unsigned( 91 , 8)),
                    2 => std_logic_vector(to_unsigned( 80 , 8)),
                    3 => std_logic_vector(to_unsigned( 105 , 8)),
                    4 => std_logic_vector(to_unsigned( 99 , 8)),
                    5 => std_logic_vector(to_unsigned( 65 , 8)),
                    6 => std_logic_vector(to_unsigned( 18 , 8)),
                    7 => std_logic_vector(to_unsigned( 48 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1041 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),
                    1 => std_logic_vector(to_unsigned( 91 , 8)),
                    2 => std_logic_vector(to_unsigned( 36 , 8)),
                    3 => std_logic_vector(to_unsigned( 23 , 8)),
                    4 => std_logic_vector(to_unsigned( 1 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 49 , 8)),
                    7 => std_logic_vector(to_unsigned( 30 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1042 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),
                    1 => std_logic_vector(to_unsigned( 91 , 8)),
                    2 => std_logic_vector(to_unsigned( 36 , 8)),
                    3 => std_logic_vector(to_unsigned( 23 , 8)),
                    4 => std_logic_vector(to_unsigned( 1 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 49 , 8)),
                    7 => std_logic_vector(to_unsigned( 30 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1043 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 2, 8)),
                    1 => std_logic_vector(to_unsigned( 50 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 122 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 32 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1044 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 10 , 8)),
                    3 => std_logic_vector(to_unsigned( 44 , 8)),
                    4 => std_logic_vector(to_unsigned( 85 , 8)),
                    5 => std_logic_vector(to_unsigned( 19 , 8)),
                    6 => std_logic_vector(to_unsigned( 48 , 8)),
                    7 => std_logic_vector(to_unsigned( 53 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1045 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 10 , 8)),
                    3 => std_logic_vector(to_unsigned( 44 , 8)),
                    4 => std_logic_vector(to_unsigned( 85 , 8)),
                    5 => std_logic_vector(to_unsigned( 19 , 8)),
                    6 => std_logic_vector(to_unsigned( 48 , 8)),
                    7 => std_logic_vector(to_unsigned( 53 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1046 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 42 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 7 , 8)),
                    4 => std_logic_vector(to_unsigned( 121 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 27 , 8)),
                    7 => std_logic_vector(to_unsigned( 113 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1047 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),
                    1 => std_logic_vector(to_unsigned( 107 , 8)),
                    2 => std_logic_vector(to_unsigned( 34 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 43 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 116 , 8)),
                    7 => std_logic_vector(to_unsigned( 20 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1048 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),
                    1 => std_logic_vector(to_unsigned( 107 , 8)),
                    2 => std_logic_vector(to_unsigned( 34 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 43 , 8)),
                    5 => std_logic_vector(to_unsigned( 96 , 8)),
                    6 => std_logic_vector(to_unsigned( 116 , 8)),
                    7 => std_logic_vector(to_unsigned( 20 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1049 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 39, 8)),
                    1 => std_logic_vector(to_unsigned( 84 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 107 , 8)),
                    4 => std_logic_vector(to_unsigned( 80 , 8)),
                    5 => std_logic_vector(to_unsigned( 18 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 31 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1050 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 118, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 78 , 8)),
                    3 => std_logic_vector(to_unsigned( 6 , 8)),
                    4 => std_logic_vector(to_unsigned( 19 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 113 , 8)),
                    7 => std_logic_vector(to_unsigned( 69 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1051 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 118, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 78 , 8)),
                    3 => std_logic_vector(to_unsigned( 6 , 8)),
                    4 => std_logic_vector(to_unsigned( 19 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 113 , 8)),
                    7 => std_logic_vector(to_unsigned( 69 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1052 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 100 , 8)),
                    2 => std_logic_vector(to_unsigned( 20 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 87 , 8)),
                    7 => std_logic_vector(to_unsigned( 29 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1053 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 5 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 34 , 8)),
                    6 => std_logic_vector(to_unsigned( 113 , 8)),
                    7 => std_logic_vector(to_unsigned( 13 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1054 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 5 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 64 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 34 , 8)),
                    6 => std_logic_vector(to_unsigned( 113 , 8)),
                    7 => std_logic_vector(to_unsigned( 13 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1055 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),
                    1 => std_logic_vector(to_unsigned( 39 , 8)),
                    2 => std_logic_vector(to_unsigned( 78 , 8)),
                    3 => std_logic_vector(to_unsigned( 63 , 8)),
                    4 => std_logic_vector(to_unsigned( 99 , 8)),
                    5 => std_logic_vector(to_unsigned( 33 , 8)),
                    6 => std_logic_vector(to_unsigned( 69 , 8)),
                    7 => std_logic_vector(to_unsigned( 21 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1056 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 86 , 8)),
                    3 => std_logic_vector(to_unsigned( 53 , 8)),
                    4 => std_logic_vector(to_unsigned( 75 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1057 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 86 , 8)),
                    3 => std_logic_vector(to_unsigned( 53 , 8)),
                    4 => std_logic_vector(to_unsigned( 75 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1058 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 2, 8)),
                    1 => std_logic_vector(to_unsigned( 98 , 8)),
                    2 => std_logic_vector(to_unsigned( 89 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 119 , 8)),
                    5 => std_logic_vector(to_unsigned( 19 , 8)),
                    6 => std_logic_vector(to_unsigned( 29 , 8)),
                    7 => std_logic_vector(to_unsigned( 7 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1059 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 80 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 105 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 29 , 8)),
                    6 => std_logic_vector(to_unsigned( 123 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1060 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 80 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 105 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 29 , 8)),
                    6 => std_logic_vector(to_unsigned( 123 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1061 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 29 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 120 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 81 , 8)),
                    7 => std_logic_vector(to_unsigned( 23 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1062 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 45, 8)),
                    1 => std_logic_vector(to_unsigned( 24 , 8)),
                    2 => std_logic_vector(to_unsigned( 83 , 8)),
                    3 => std_logic_vector(to_unsigned( 112 , 8)),
                    4 => std_logic_vector(to_unsigned( 72 , 8)),
                    5 => std_logic_vector(to_unsigned( 41 , 8)),
                    6 => std_logic_vector(to_unsigned( 76 , 8)),
                    7 => std_logic_vector(to_unsigned( 120 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1063 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 45, 8)),
                    1 => std_logic_vector(to_unsigned( 24 , 8)),
                    2 => std_logic_vector(to_unsigned( 83 , 8)),
                    3 => std_logic_vector(to_unsigned( 112 , 8)),
                    4 => std_logic_vector(to_unsigned( 72 , 8)),
                    5 => std_logic_vector(to_unsigned( 41 , 8)),
                    6 => std_logic_vector(to_unsigned( 76 , 8)),
                    7 => std_logic_vector(to_unsigned( 120 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1064 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 43 , 8)),
                    3 => std_logic_vector(to_unsigned( 65 , 8)),
                    4 => std_logic_vector(to_unsigned( 38 , 8)),
                    5 => std_logic_vector(to_unsigned( 61 , 8)),
                    6 => std_logic_vector(to_unsigned( 16 , 8)),
                    7 => std_logic_vector(to_unsigned( 88 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1065 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 35 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 122 , 8)),
                    4 => std_logic_vector(to_unsigned( 49 , 8)),
                    5 => std_logic_vector(to_unsigned( 30 , 8)),
                    6 => std_logic_vector(to_unsigned( 20 , 8)),
                    7 => std_logic_vector(to_unsigned( 96 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1066 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 35 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 122 , 8)),
                    4 => std_logic_vector(to_unsigned( 49 , 8)),
                    5 => std_logic_vector(to_unsigned( 30 , 8)),
                    6 => std_logic_vector(to_unsigned( 20 , 8)),
                    7 => std_logic_vector(to_unsigned( 96 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1067 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 17, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 51 , 8)),
                    3 => std_logic_vector(to_unsigned( 75 , 8)),
                    4 => std_logic_vector(to_unsigned( 60 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 83 , 8)),
                    7 => std_logic_vector(to_unsigned( 25 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1068 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 112, 8)),
                    1 => std_logic_vector(to_unsigned( 124 , 8)),
                    2 => std_logic_vector(to_unsigned( 54 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 63 , 8)),
                    5 => std_logic_vector(to_unsigned( 38 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 98 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1069 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 112, 8)),
                    1 => std_logic_vector(to_unsigned( 124 , 8)),
                    2 => std_logic_vector(to_unsigned( 54 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 63 , 8)),
                    5 => std_logic_vector(to_unsigned( 38 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 98 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1070 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 20 , 8)),
                    3 => std_logic_vector(to_unsigned( 10 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 55 , 8)),
                    6 => std_logic_vector(to_unsigned( 102 , 8)),
                    7 => std_logic_vector(to_unsigned( 98 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1071 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),
                    1 => std_logic_vector(to_unsigned( 117 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 79 , 8)),
                    4 => std_logic_vector(to_unsigned( 13 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 99 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1072 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),
                    1 => std_logic_vector(to_unsigned( 117 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 79 , 8)),
                    4 => std_logic_vector(to_unsigned( 13 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 99 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1073 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 66 , 8)),
                    2 => std_logic_vector(to_unsigned( 116 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 19 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 89 , 8)),
                    7 => std_logic_vector(to_unsigned( 46 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1074 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 82, 8)),
                    1 => std_logic_vector(to_unsigned( 44 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 103 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 20 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1075 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 82, 8)),
                    1 => std_logic_vector(to_unsigned( 44 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 103 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 20 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1076 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 110, 8)),
                    1 => std_logic_vector(to_unsigned( 17 , 8)),
                    2 => std_logic_vector(to_unsigned( 83 , 8)),
                    3 => std_logic_vector(to_unsigned( 27 , 8)),
                    4 => std_logic_vector(to_unsigned( 77 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 70 , 8)),
                    7 => std_logic_vector(to_unsigned( 5 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1077 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 112 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 31 , 8)),
                    4 => std_logic_vector(to_unsigned( 85 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 81 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1078 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 112 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 31 , 8)),
                    4 => std_logic_vector(to_unsigned( 85 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 81 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1079 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 109, 8)),
                    1 => std_logic_vector(to_unsigned( 86 , 8)),
                    2 => std_logic_vector(to_unsigned( 20 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 113 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1080 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),
                    1 => std_logic_vector(to_unsigned( 85 , 8)),
                    2 => std_logic_vector(to_unsigned( 48 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 124 , 8)),
                    6 => std_logic_vector(to_unsigned( 111 , 8)),
                    7 => std_logic_vector(to_unsigned( 81 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1081 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),
                    1 => std_logic_vector(to_unsigned( 85 , 8)),
                    2 => std_logic_vector(to_unsigned( 48 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 124 , 8)),
                    6 => std_logic_vector(to_unsigned( 111 , 8)),
                    7 => std_logic_vector(to_unsigned( 81 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1082 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 117 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 1 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 56 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1083 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),
                    1 => std_logic_vector(to_unsigned( 50 , 8)),
                    2 => std_logic_vector(to_unsigned( 84 , 8)),
                    3 => std_logic_vector(to_unsigned( 27 , 8)),
                    4 => std_logic_vector(to_unsigned( 42 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 121 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1084 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),
                    1 => std_logic_vector(to_unsigned( 50 , 8)),
                    2 => std_logic_vector(to_unsigned( 84 , 8)),
                    3 => std_logic_vector(to_unsigned( 27 , 8)),
                    4 => std_logic_vector(to_unsigned( 42 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 121 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1085 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),
                    1 => std_logic_vector(to_unsigned( 94 , 8)),
                    2 => std_logic_vector(to_unsigned( 70 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 121 , 8)),
                    5 => std_logic_vector(to_unsigned( 22 , 8)),
                    6 => std_logic_vector(to_unsigned( 65 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1086 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 117 , 8)),
                    2 => std_logic_vector(to_unsigned( 108 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 86 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 4 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1087 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 117 , 8)),
                    2 => std_logic_vector(to_unsigned( 108 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 86 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 4 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1088 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 43 , 8)),
                    3 => std_logic_vector(to_unsigned( 17 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 35 , 8)),
                    7 => std_logic_vector(to_unsigned( 117 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1089 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),
                    1 => std_logic_vector(to_unsigned( 110 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 15 , 8)),
                    4 => std_logic_vector(to_unsigned( 76 , 8)),
                    5 => std_logic_vector(to_unsigned( 30 , 8)),
                    6 => std_logic_vector(to_unsigned( 58 , 8)),
                    7 => std_logic_vector(to_unsigned( 10 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1090 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),
                    1 => std_logic_vector(to_unsigned( 110 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 15 , 8)),
                    4 => std_logic_vector(to_unsigned( 76 , 8)),
                    5 => std_logic_vector(to_unsigned( 30 , 8)),
                    6 => std_logic_vector(to_unsigned( 58 , 8)),
                    7 => std_logic_vector(to_unsigned( 10 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1091 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 65, 8)),
                    1 => std_logic_vector(to_unsigned( 72 , 8)),
                    2 => std_logic_vector(to_unsigned( 85 , 8)),
                    3 => std_logic_vector(to_unsigned( 108 , 8)),
                    4 => std_logic_vector(to_unsigned( 14 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 29 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1092 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),
                    1 => std_logic_vector(to_unsigned( 54 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 4 , 8)),
                    5 => std_logic_vector(to_unsigned( 112 , 8)),
                    6 => std_logic_vector(to_unsigned( 68 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1093 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),
                    1 => std_logic_vector(to_unsigned( 54 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 4 , 8)),
                    5 => std_logic_vector(to_unsigned( 112 , 8)),
                    6 => std_logic_vector(to_unsigned( 68 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1094 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),
                    1 => std_logic_vector(to_unsigned( 40 , 8)),
                    2 => std_logic_vector(to_unsigned( 102 , 8)),
                    3 => std_logic_vector(to_unsigned( 57 , 8)),
                    4 => std_logic_vector(to_unsigned( 64 , 8)),
                    5 => std_logic_vector(to_unsigned( 32 , 8)),
                    6 => std_logic_vector(to_unsigned( 21 , 8)),
                    7 => std_logic_vector(to_unsigned( 92 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1095 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 25 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 46 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1096 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 25 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 46 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1097 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 75 , 8)),
                    3 => std_logic_vector(to_unsigned( 120 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 88 , 8)),
                    7 => std_logic_vector(to_unsigned( 25 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1098 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),
                    1 => std_logic_vector(to_unsigned( 81 , 8)),
                    2 => std_logic_vector(to_unsigned( 9 , 8)),
                    3 => std_logic_vector(to_unsigned( 117 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 29 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1099 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),
                    1 => std_logic_vector(to_unsigned( 81 , 8)),
                    2 => std_logic_vector(to_unsigned( 9 , 8)),
                    3 => std_logic_vector(to_unsigned( 117 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 29 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1100 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 97, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 54 , 8)),
                    3 => std_logic_vector(to_unsigned( 25 , 8)),
                    4 => std_logic_vector(to_unsigned( 18 , 8)),
                    5 => std_logic_vector(to_unsigned( 103 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 90 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1101 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),
                    1 => std_logic_vector(to_unsigned( 99 , 8)),
                    2 => std_logic_vector(to_unsigned( 12 , 8)),
                    3 => std_logic_vector(to_unsigned( 121 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 76 , 8)),
                    6 => std_logic_vector(to_unsigned( 41 , 8)),
                    7 => std_logic_vector(to_unsigned( 64 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1102 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),
                    1 => std_logic_vector(to_unsigned( 99 , 8)),
                    2 => std_logic_vector(to_unsigned( 12 , 8)),
                    3 => std_logic_vector(to_unsigned( 121 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 76 , 8)),
                    6 => std_logic_vector(to_unsigned( 41 , 8)),
                    7 => std_logic_vector(to_unsigned( 64 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1103 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),
                    1 => std_logic_vector(to_unsigned( 76 , 8)),
                    2 => std_logic_vector(to_unsigned( 109 , 8)),
                    3 => std_logic_vector(to_unsigned( 44 , 8)),
                    4 => std_logic_vector(to_unsigned( 94 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 90 , 8)),
                    7 => std_logic_vector(to_unsigned( 3 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1104 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),
                    1 => std_logic_vector(to_unsigned( 95 , 8)),
                    2 => std_logic_vector(to_unsigned( 52 , 8)),
                    3 => std_logic_vector(to_unsigned( 19 , 8)),
                    4 => std_logic_vector(to_unsigned( 108 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 85 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1105 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),
                    1 => std_logic_vector(to_unsigned( 95 , 8)),
                    2 => std_logic_vector(to_unsigned( 52 , 8)),
                    3 => std_logic_vector(to_unsigned( 19 , 8)),
                    4 => std_logic_vector(to_unsigned( 108 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 85 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1106 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 38, 8)),
                    1 => std_logic_vector(to_unsigned( 110 , 8)),
                    2 => std_logic_vector(to_unsigned( 61 , 8)),
                    3 => std_logic_vector(to_unsigned( 77 , 8)),
                    4 => std_logic_vector(to_unsigned( 17 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 118 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1107 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 2 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 77 , 8)),
                    5 => std_logic_vector(to_unsigned( 39 , 8)),
                    6 => std_logic_vector(to_unsigned( 106 , 8)),
                    7 => std_logic_vector(to_unsigned( 29 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1108 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 2 , 8)),
                    3 => std_logic_vector(to_unsigned( 87 , 8)),
                    4 => std_logic_vector(to_unsigned( 77 , 8)),
                    5 => std_logic_vector(to_unsigned( 39 , 8)),
                    6 => std_logic_vector(to_unsigned( 106 , 8)),
                    7 => std_logic_vector(to_unsigned( 29 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1109 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),
                    1 => std_logic_vector(to_unsigned( 17 , 8)),
                    2 => std_logic_vector(to_unsigned( 116 , 8)),
                    3 => std_logic_vector(to_unsigned( 60 , 8)),
                    4 => std_logic_vector(to_unsigned( 24 , 8)),
                    5 => std_logic_vector(to_unsigned( 42 , 8)),
                    6 => std_logic_vector(to_unsigned( 68 , 8)),
                    7 => std_logic_vector(to_unsigned( 81 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1110 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),
                    1 => std_logic_vector(to_unsigned( 112 , 8)),
                    2 => std_logic_vector(to_unsigned( 49 , 8)),
                    3 => std_logic_vector(to_unsigned( 75 , 8)),
                    4 => std_logic_vector(to_unsigned( 40 , 8)),
                    5 => std_logic_vector(to_unsigned( 116 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1111 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),
                    1 => std_logic_vector(to_unsigned( 112 , 8)),
                    2 => std_logic_vector(to_unsigned( 49 , 8)),
                    3 => std_logic_vector(to_unsigned( 75 , 8)),
                    4 => std_logic_vector(to_unsigned( 40 , 8)),
                    5 => std_logic_vector(to_unsigned( 116 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1112 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 51, 8)),
                    1 => std_logic_vector(to_unsigned( 38 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 123 , 8)),
                    4 => std_logic_vector(to_unsigned( 11 , 8)),
                    5 => std_logic_vector(to_unsigned( 17 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 112 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1113 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 2, 8)),
                    1 => std_logic_vector(to_unsigned( 66 , 8)),
                    2 => std_logic_vector(to_unsigned( 99 , 8)),
                    3 => std_logic_vector(to_unsigned( 89 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 74 , 8)),
                    6 => std_logic_vector(to_unsigned( 57 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1114 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 2, 8)),
                    1 => std_logic_vector(to_unsigned( 66 , 8)),
                    2 => std_logic_vector(to_unsigned( 99 , 8)),
                    3 => std_logic_vector(to_unsigned( 89 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 74 , 8)),
                    6 => std_logic_vector(to_unsigned( 57 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1115 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 40, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 21 , 8)),
                    3 => std_logic_vector(to_unsigned( 16 , 8)),
                    4 => std_logic_vector(to_unsigned( 9 , 8)),
                    5 => std_logic_vector(to_unsigned( 28 , 8)),
                    6 => std_logic_vector(to_unsigned( 90 , 8)),
                    7 => std_logic_vector(to_unsigned( 121 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1116 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),
                    1 => std_logic_vector(to_unsigned( 33 , 8)),
                    2 => std_logic_vector(to_unsigned( 79 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 93 , 8)),
                    7 => std_logic_vector(to_unsigned( 27 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1117 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),
                    1 => std_logic_vector(to_unsigned( 33 , 8)),
                    2 => std_logic_vector(to_unsigned( 79 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 93 , 8)),
                    7 => std_logic_vector(to_unsigned( 27 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1118 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),
                    1 => std_logic_vector(to_unsigned( 19 , 8)),
                    2 => std_logic_vector(to_unsigned( 100 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 119 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 82 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1119 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 97, 8)),
                    1 => std_logic_vector(to_unsigned( 60 , 8)),
                    2 => std_logic_vector(to_unsigned( 114 , 8)),
                    3 => std_logic_vector(to_unsigned( 56 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 102 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 46 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1120 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 97, 8)),
                    1 => std_logic_vector(to_unsigned( 60 , 8)),
                    2 => std_logic_vector(to_unsigned( 114 , 8)),
                    3 => std_logic_vector(to_unsigned( 56 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 102 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 46 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1121 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 86 , 8)),
                    4 => std_logic_vector(to_unsigned( 13 , 8)),
                    5 => std_logic_vector(to_unsigned( 22 , 8)),
                    6 => std_logic_vector(to_unsigned( 35 , 8)),
                    7 => std_logic_vector(to_unsigned( 9 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1122 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 100 , 8)),
                    3 => std_logic_vector(to_unsigned( 104 , 8)),
                    4 => std_logic_vector(to_unsigned( 24 , 8)),
                    5 => std_logic_vector(to_unsigned( 32 , 8)),
                    6 => std_logic_vector(to_unsigned( 74 , 8)),
                    7 => std_logic_vector(to_unsigned( 121 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1123 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 100 , 8)),
                    3 => std_logic_vector(to_unsigned( 104 , 8)),
                    4 => std_logic_vector(to_unsigned( 24 , 8)),
                    5 => std_logic_vector(to_unsigned( 32 , 8)),
                    6 => std_logic_vector(to_unsigned( 74 , 8)),
                    7 => std_logic_vector(to_unsigned( 121 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1124 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),
                    1 => std_logic_vector(to_unsigned( 111 , 8)),
                    2 => std_logic_vector(to_unsigned( 2 , 8)),
                    3 => std_logic_vector(to_unsigned( 69 , 8)),
                    4 => std_logic_vector(to_unsigned( 41 , 8)),
                    5 => std_logic_vector(to_unsigned( 103 , 8)),
                    6 => std_logic_vector(to_unsigned( 90 , 8)),
                    7 => std_logic_vector(to_unsigned( 115 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1125 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 21 , 8)),
                    2 => std_logic_vector(to_unsigned( 12 , 8)),
                    3 => std_logic_vector(to_unsigned( 73 , 8)),
                    4 => std_logic_vector(to_unsigned( 31 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 109 , 8)),
                    7 => std_logic_vector(to_unsigned( 8 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1126 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 21 , 8)),
                    2 => std_logic_vector(to_unsigned( 12 , 8)),
                    3 => std_logic_vector(to_unsigned( 73 , 8)),
                    4 => std_logic_vector(to_unsigned( 31 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 109 , 8)),
                    7 => std_logic_vector(to_unsigned( 8 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1127 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 25, 8)),
                    1 => std_logic_vector(to_unsigned( 94 , 8)),
                    2 => std_logic_vector(to_unsigned( 62 , 8)),
                    3 => std_logic_vector(to_unsigned( 39 , 8)),
                    4 => std_logic_vector(to_unsigned( 7 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 18 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1128 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),
                    1 => std_logic_vector(to_unsigned( 85 , 8)),
                    2 => std_logic_vector(to_unsigned( 40 , 8)),
                    3 => std_logic_vector(to_unsigned( 108 , 8)),
                    4 => std_logic_vector(to_unsigned( 115 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 94 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1129 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),
                    1 => std_logic_vector(to_unsigned( 85 , 8)),
                    2 => std_logic_vector(to_unsigned( 40 , 8)),
                    3 => std_logic_vector(to_unsigned( 108 , 8)),
                    4 => std_logic_vector(to_unsigned( 115 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 94 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1130 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),
                    1 => std_logic_vector(to_unsigned( 6 , 8)),
                    2 => std_logic_vector(to_unsigned( 15 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 70 , 8)),
                    5 => std_logic_vector(to_unsigned( 92 , 8)),
                    6 => std_logic_vector(to_unsigned( 54 , 8)),
                    7 => std_logic_vector(to_unsigned( 46 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1131 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 91 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 109 , 8)),
                    4 => std_logic_vector(to_unsigned( 123 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 38 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1132 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 91 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 109 , 8)),
                    4 => std_logic_vector(to_unsigned( 123 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 38 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1133 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 29 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 68 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 101 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1134 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 99, 8)),
                    1 => std_logic_vector(to_unsigned( 7 , 8)),
                    2 => std_logic_vector(to_unsigned( 60 , 8)),
                    3 => std_logic_vector(to_unsigned( 111 , 8)),
                    4 => std_logic_vector(to_unsigned( 76 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 44 , 8)),
                    7 => std_logic_vector(to_unsigned( 18 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1135 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 99, 8)),
                    1 => std_logic_vector(to_unsigned( 7 , 8)),
                    2 => std_logic_vector(to_unsigned( 60 , 8)),
                    3 => std_logic_vector(to_unsigned( 111 , 8)),
                    4 => std_logic_vector(to_unsigned( 76 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 44 , 8)),
                    7 => std_logic_vector(to_unsigned( 18 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1136 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),
                    1 => std_logic_vector(to_unsigned( 120 , 8)),
                    2 => std_logic_vector(to_unsigned( 46 , 8)),
                    3 => std_logic_vector(to_unsigned( 10 , 8)),
                    4 => std_logic_vector(to_unsigned( 23 , 8)),
                    5 => std_logic_vector(to_unsigned( 37 , 8)),
                    6 => std_logic_vector(to_unsigned( 90 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1137 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 13 , 8)),
                    3 => std_logic_vector(to_unsigned( 103 , 8)),
                    4 => std_logic_vector(to_unsigned( 23 , 8)),
                    5 => std_logic_vector(to_unsigned( 17 , 8)),
                    6 => std_logic_vector(to_unsigned( 112 , 8)),
                    7 => std_logic_vector(to_unsigned( 61 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1138 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 13 , 8)),
                    3 => std_logic_vector(to_unsigned( 103 , 8)),
                    4 => std_logic_vector(to_unsigned( 23 , 8)),
                    5 => std_logic_vector(to_unsigned( 17 , 8)),
                    6 => std_logic_vector(to_unsigned( 112 , 8)),
                    7 => std_logic_vector(to_unsigned( 61 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1139 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),
                    1 => std_logic_vector(to_unsigned( 19 , 8)),
                    2 => std_logic_vector(to_unsigned( 24 , 8)),
                    3 => std_logic_vector(to_unsigned( 49 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 61 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1140 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 15 , 8)),
                    3 => std_logic_vector(to_unsigned( 110 , 8)),
                    4 => std_logic_vector(to_unsigned( 32 , 8)),
                    5 => std_logic_vector(to_unsigned( 70 , 8)),
                    6 => std_logic_vector(to_unsigned( 60 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1141 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 15 , 8)),
                    3 => std_logic_vector(to_unsigned( 110 , 8)),
                    4 => std_logic_vector(to_unsigned( 32 , 8)),
                    5 => std_logic_vector(to_unsigned( 70 , 8)),
                    6 => std_logic_vector(to_unsigned( 60 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1142 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 68 , 8)),
                    2 => std_logic_vector(to_unsigned( 39 , 8)),
                    3 => std_logic_vector(to_unsigned( 81 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 72 , 8)),
                    6 => std_logic_vector(to_unsigned( 22 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1143 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 108 , 8)),
                    4 => std_logic_vector(to_unsigned( 53 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 26 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1144 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 108 , 8)),
                    4 => std_logic_vector(to_unsigned( 53 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 26 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1145 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 102 , 8)),
                    3 => std_logic_vector(to_unsigned( 63 , 8)),
                    4 => std_logic_vector(to_unsigned( 124 , 8)),
                    5 => std_logic_vector(to_unsigned( 17 , 8)),
                    6 => std_logic_vector(to_unsigned( 25 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1146 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 85 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 112 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1147 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 85 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 112 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1148 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 23 , 8)),
                    4 => std_logic_vector(to_unsigned( 73 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 27 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1149 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),
                    1 => std_logic_vector(to_unsigned( 72 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 111 , 8)),
                    4 => std_logic_vector(to_unsigned( 23 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 54 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1150 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),
                    1 => std_logic_vector(to_unsigned( 72 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 111 , 8)),
                    4 => std_logic_vector(to_unsigned( 23 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 54 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1151 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),
                    1 => std_logic_vector(to_unsigned( 119 , 8)),
                    2 => std_logic_vector(to_unsigned( 39 , 8)),
                    3 => std_logic_vector(to_unsigned( 17 , 8)),
                    4 => std_logic_vector(to_unsigned( 86 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 59 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1152 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 48 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 66 , 8)),
                    5 => std_logic_vector(to_unsigned( 56 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 111 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1153 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 48 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 66 , 8)),
                    5 => std_logic_vector(to_unsigned( 56 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 111 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1154 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 64 , 8)),
                    3 => std_logic_vector(to_unsigned( 44 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 84 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 56 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1155 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 2 , 8)),
                    3 => std_logic_vector(to_unsigned( 91 , 8)),
                    4 => std_logic_vector(to_unsigned( 69 , 8)),
                    5 => std_logic_vector(to_unsigned( 19 , 8)),
                    6 => std_logic_vector(to_unsigned( 23 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1156 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 2 , 8)),
                    3 => std_logic_vector(to_unsigned( 91 , 8)),
                    4 => std_logic_vector(to_unsigned( 69 , 8)),
                    5 => std_logic_vector(to_unsigned( 19 , 8)),
                    6 => std_logic_vector(to_unsigned( 23 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1157 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 46 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 85 , 8)),
                    4 => std_logic_vector(to_unsigned( 34 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 30 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1158 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 40 , 8)),
                    3 => std_logic_vector(to_unsigned( 113 , 8)),
                    4 => std_logic_vector(to_unsigned( 54 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 46 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1159 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 40 , 8)),
                    3 => std_logic_vector(to_unsigned( 113 , 8)),
                    4 => std_logic_vector(to_unsigned( 54 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 46 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1160 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),
                    1 => std_logic_vector(to_unsigned( 27 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 118 , 8)),
                    5 => std_logic_vector(to_unsigned( 65 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 69 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1161 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),
                    1 => std_logic_vector(to_unsigned( 108 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 42 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1162 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),
                    1 => std_logic_vector(to_unsigned( 108 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 42 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1163 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 19 , 8)),
                    2 => std_logic_vector(to_unsigned( 58 , 8)),
                    3 => std_logic_vector(to_unsigned( 93 , 8)),
                    4 => std_logic_vector(to_unsigned( 66 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 115 , 8)),
                    7 => std_logic_vector(to_unsigned( 43 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1164 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 15 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 101 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 45 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1165 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 15 , 8)),
                    2 => std_logic_vector(to_unsigned( 25 , 8)),
                    3 => std_logic_vector(to_unsigned( 101 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 45 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1166 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 67, 8)),
                    1 => std_logic_vector(to_unsigned( 54 , 8)),
                    2 => std_logic_vector(to_unsigned( 113 , 8)),
                    3 => std_logic_vector(to_unsigned( 60 , 8)),
                    4 => std_logic_vector(to_unsigned( 83 , 8)),
                    5 => std_logic_vector(to_unsigned( 46 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1167 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 105, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 26 , 8)),
                    3 => std_logic_vector(to_unsigned( 53 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 57 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1168 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 105, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 26 , 8)),
                    3 => std_logic_vector(to_unsigned( 53 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 57 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1169 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),
                    1 => std_logic_vector(to_unsigned( 119 , 8)),
                    2 => std_logic_vector(to_unsigned( 47 , 8)),
                    3 => std_logic_vector(to_unsigned( 100 , 8)),
                    4 => std_logic_vector(to_unsigned( 53 , 8)),
                    5 => std_logic_vector(to_unsigned( 0 , 8)),
                    6 => std_logic_vector(to_unsigned( 105 , 8)),
                    7 => std_logic_vector(to_unsigned( 39 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1170 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),
                    1 => std_logic_vector(to_unsigned( 79 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 29 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 3 , 8)),
                    7 => std_logic_vector(to_unsigned( 22 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1171 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),
                    1 => std_logic_vector(to_unsigned( 79 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 29 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 3 , 8)),
                    7 => std_logic_vector(to_unsigned( 22 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1172 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),
                    1 => std_logic_vector(to_unsigned( 29 , 8)),
                    2 => std_logic_vector(to_unsigned( 65 , 8)),
                    3 => std_logic_vector(to_unsigned( 88 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 102 , 8)),
                    6 => std_logic_vector(to_unsigned( 44 , 8)),
                    7 => std_logic_vector(to_unsigned( 1 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1173 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 45, 8)),
                    1 => std_logic_vector(to_unsigned( 54 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 120 , 8)),
                    4 => std_logic_vector(to_unsigned( 69 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1174 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 45, 8)),
                    1 => std_logic_vector(to_unsigned( 54 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 120 , 8)),
                    4 => std_logic_vector(to_unsigned( 69 , 8)),
                    5 => std_logic_vector(to_unsigned( 4 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1175 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 9, 8)),
                    1 => std_logic_vector(to_unsigned( 95 , 8)),
                    2 => std_logic_vector(to_unsigned( 78 , 8)),
                    3 => std_logic_vector(to_unsigned( 43 , 8)),
                    4 => std_logic_vector(to_unsigned( 34 , 8)),
                    5 => std_logic_vector(to_unsigned( 23 , 8)),
                    6 => std_logic_vector(to_unsigned( 107 , 8)),
                    7 => std_logic_vector(to_unsigned( 57 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1176 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),
                    1 => std_logic_vector(to_unsigned( 0 , 8)),
                    2 => std_logic_vector(to_unsigned( 80 , 8)),
                    3 => std_logic_vector(to_unsigned( 75 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 14 , 8)),
                    6 => std_logic_vector(to_unsigned( 91 , 8)),
                    7 => std_logic_vector(to_unsigned( 71 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1177 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),
                    1 => std_logic_vector(to_unsigned( 0 , 8)),
                    2 => std_logic_vector(to_unsigned( 80 , 8)),
                    3 => std_logic_vector(to_unsigned( 75 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 14 , 8)),
                    6 => std_logic_vector(to_unsigned( 91 , 8)),
                    7 => std_logic_vector(to_unsigned( 71 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1178 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 76, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 64 , 8)),
                    3 => std_logic_vector(to_unsigned( 124 , 8)),
                    4 => std_logic_vector(to_unsigned( 97 , 8)),
                    5 => std_logic_vector(to_unsigned( 115 , 8)),
                    6 => std_logic_vector(to_unsigned( 16 , 8)),
                    7 => std_logic_vector(to_unsigned( 57 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1179 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),
                    1 => std_logic_vector(to_unsigned( 64 , 8)),
                    2 => std_logic_vector(to_unsigned( 54 , 8)),
                    3 => std_logic_vector(to_unsigned( 17 , 8)),
                    4 => std_logic_vector(to_unsigned( 11 , 8)),
                    5 => std_logic_vector(to_unsigned( 74 , 8)),
                    6 => std_logic_vector(to_unsigned( 1 , 8)),
                    7 => std_logic_vector(to_unsigned( 121 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1180 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),
                    1 => std_logic_vector(to_unsigned( 64 , 8)),
                    2 => std_logic_vector(to_unsigned( 54 , 8)),
                    3 => std_logic_vector(to_unsigned( 17 , 8)),
                    4 => std_logic_vector(to_unsigned( 11 , 8)),
                    5 => std_logic_vector(to_unsigned( 74 , 8)),
                    6 => std_logic_vector(to_unsigned( 1 , 8)),
                    7 => std_logic_vector(to_unsigned( 121 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1181 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 41, 8)),
                    1 => std_logic_vector(to_unsigned( 71 , 8)),
                    2 => std_logic_vector(to_unsigned( 12 , 8)),
                    3 => std_logic_vector(to_unsigned( 45 , 8)),
                    4 => std_logic_vector(to_unsigned( 124 , 8)),
                    5 => std_logic_vector(to_unsigned( 23 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 96 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1182 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 104 , 8)),
                    3 => std_logic_vector(to_unsigned( 79 , 8)),
                    4 => std_logic_vector(to_unsigned( 122 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 64 , 8)),
                    7 => std_logic_vector(to_unsigned( 5 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1183 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 104 , 8)),
                    3 => std_logic_vector(to_unsigned( 79 , 8)),
                    4 => std_logic_vector(to_unsigned( 122 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 64 , 8)),
                    7 => std_logic_vector(to_unsigned( 5 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1184 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 66 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 41 , 8)),
                    4 => std_logic_vector(to_unsigned( 91 , 8)),
                    5 => std_logic_vector(to_unsigned( 112 , 8)),
                    6 => std_logic_vector(to_unsigned( 48 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1185 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),
                    1 => std_logic_vector(to_unsigned( 82 , 8)),
                    2 => std_logic_vector(to_unsigned( 50 , 8)),
                    3 => std_logic_vector(to_unsigned( 97 , 8)),
                    4 => std_logic_vector(to_unsigned( 68 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 102 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1186 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),
                    1 => std_logic_vector(to_unsigned( 82 , 8)),
                    2 => std_logic_vector(to_unsigned( 50 , 8)),
                    3 => std_logic_vector(to_unsigned( 97 , 8)),
                    4 => std_logic_vector(to_unsigned( 68 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 102 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1187 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),
                    1 => std_logic_vector(to_unsigned( 111 , 8)),
                    2 => std_logic_vector(to_unsigned( 19 , 8)),
                    3 => std_logic_vector(to_unsigned( 123 , 8)),
                    4 => std_logic_vector(to_unsigned( 13 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 106 , 8)),
                    7 => std_logic_vector(to_unsigned( 74 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1188 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),
                    1 => std_logic_vector(to_unsigned( 72 , 8)),
                    2 => std_logic_vector(to_unsigned( 68 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 27 , 8)),
                    5 => std_logic_vector(to_unsigned( 8 , 8)),
                    6 => std_logic_vector(to_unsigned( 15 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1189 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),
                    1 => std_logic_vector(to_unsigned( 72 , 8)),
                    2 => std_logic_vector(to_unsigned( 68 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 27 , 8)),
                    5 => std_logic_vector(to_unsigned( 8 , 8)),
                    6 => std_logic_vector(to_unsigned( 15 , 8)),
                    7 => std_logic_vector(to_unsigned( 114 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1190 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 85 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 81 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 51 , 8)),
                    6 => std_logic_vector(to_unsigned( 28 , 8)),
                    7 => std_logic_vector(to_unsigned( 1 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1191 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 76 , 8)),
                    4 => std_logic_vector(to_unsigned( 68 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 116 , 8)),
                    7 => std_logic_vector(to_unsigned( 47 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1192 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 76 , 8)),
                    4 => std_logic_vector(to_unsigned( 68 , 8)),
                    5 => std_logic_vector(to_unsigned( 59 , 8)),
                    6 => std_logic_vector(to_unsigned( 116 , 8)),
                    7 => std_logic_vector(to_unsigned( 47 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1193 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 12, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 37 , 8)),
                    5 => std_logic_vector(to_unsigned( 49 , 8)),
                    6 => std_logic_vector(to_unsigned( 117 , 8)),
                    7 => std_logic_vector(to_unsigned( 7 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1194 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 12, 8)),
                    1 => std_logic_vector(to_unsigned( 90 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 86 , 8)),
                    4 => std_logic_vector(to_unsigned( 18 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 68 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1195 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 12, 8)),
                    1 => std_logic_vector(to_unsigned( 90 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 86 , 8)),
                    4 => std_logic_vector(to_unsigned( 18 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 68 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1196 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),
                    1 => std_logic_vector(to_unsigned( 119 , 8)),
                    2 => std_logic_vector(to_unsigned( 13 , 8)),
                    3 => std_logic_vector(to_unsigned( 103 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 73 , 8)),
                    6 => std_logic_vector(to_unsigned( 52 , 8)),
                    7 => std_logic_vector(to_unsigned( 19 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1197 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 9, 8)),
                    1 => std_logic_vector(to_unsigned( 101 , 8)),
                    2 => std_logic_vector(to_unsigned( 61 , 8)),
                    3 => std_logic_vector(to_unsigned( 76 , 8)),
                    4 => std_logic_vector(to_unsigned( 110 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 114 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1198 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 9, 8)),
                    1 => std_logic_vector(to_unsigned( 101 , 8)),
                    2 => std_logic_vector(to_unsigned( 61 , 8)),
                    3 => std_logic_vector(to_unsigned( 76 , 8)),
                    4 => std_logic_vector(to_unsigned( 110 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 114 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1199 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),
                    1 => std_logic_vector(to_unsigned( 34 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 114 , 8)),
                    4 => std_logic_vector(to_unsigned( 76 , 8)),
                    5 => std_logic_vector(to_unsigned( 30 , 8)),
                    6 => std_logic_vector(to_unsigned( 12 , 8)),
                    7 => std_logic_vector(to_unsigned( 42 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1200 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 82, 8)),
                    1 => std_logic_vector(to_unsigned( 6 , 8)),
                    2 => std_logic_vector(to_unsigned( 112 , 8)),
                    3 => std_logic_vector(to_unsigned( 89 , 8)),
                    4 => std_logic_vector(to_unsigned( 20 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 70 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1201 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 82, 8)),
                    1 => std_logic_vector(to_unsigned( 6 , 8)),
                    2 => std_logic_vector(to_unsigned( 112 , 8)),
                    3 => std_logic_vector(to_unsigned( 89 , 8)),
                    4 => std_logic_vector(to_unsigned( 20 , 8)),
                    5 => std_logic_vector(to_unsigned( 53 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 70 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1202 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 4, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 84 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 49 , 8)),
                    5 => std_logic_vector(to_unsigned( 24 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 61 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1203 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 80 , 8)),
                    2 => std_logic_vector(to_unsigned( 28 , 8)),
                    3 => std_logic_vector(to_unsigned( 37 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 87 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 98 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1204 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 80 , 8)),
                    2 => std_logic_vector(to_unsigned( 28 , 8)),
                    3 => std_logic_vector(to_unsigned( 37 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 87 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 98 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1205 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),
                    1 => std_logic_vector(to_unsigned( 0 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 120 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 93 , 8)),
                    7 => std_logic_vector(to_unsigned( 23 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1206 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 31 , 8)),
                    4 => std_logic_vector(to_unsigned( 22 , 8)),
                    5 => std_logic_vector(to_unsigned( 82 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1207 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 31 , 8)),
                    4 => std_logic_vector(to_unsigned( 22 , 8)),
                    5 => std_logic_vector(to_unsigned( 82 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1208 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),
                    1 => std_logic_vector(to_unsigned( 5 , 8)),
                    2 => std_logic_vector(to_unsigned( 18 , 8)),
                    3 => std_logic_vector(to_unsigned( 55 , 8)),
                    4 => std_logic_vector(to_unsigned( 98 , 8)),
                    5 => std_logic_vector(to_unsigned( 61 , 8)),
                    6 => std_logic_vector(to_unsigned( 89 , 8)),
                    7 => std_logic_vector(to_unsigned( 107 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1209 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 12, 8)),
                    1 => std_logic_vector(to_unsigned( 50 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 71 , 8)),
                    4 => std_logic_vector(to_unsigned( 18 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1210 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 12, 8)),
                    1 => std_logic_vector(to_unsigned( 50 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 71 , 8)),
                    4 => std_logic_vector(to_unsigned( 18 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1211 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),
                    1 => std_logic_vector(to_unsigned( 85 , 8)),
                    2 => std_logic_vector(to_unsigned( 35 , 8)),
                    3 => std_logic_vector(to_unsigned( 23 , 8)),
                    4 => std_logic_vector(to_unsigned( 5 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 120 , 8)),
                    7 => std_logic_vector(to_unsigned( 56 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1212 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 24 , 8)),
                    2 => std_logic_vector(to_unsigned( 52 , 8)),
                    3 => std_logic_vector(to_unsigned( 66 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 36 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 79 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1213 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),
                    1 => std_logic_vector(to_unsigned( 24 , 8)),
                    2 => std_logic_vector(to_unsigned( 52 , 8)),
                    3 => std_logic_vector(to_unsigned( 66 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 36 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 79 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1214 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),
                    1 => std_logic_vector(to_unsigned( 67 , 8)),
                    2 => std_logic_vector(to_unsigned( 101 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 8 , 8)),
                    5 => std_logic_vector(to_unsigned( 105 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1215 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 72, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 18 , 8)),
                    4 => std_logic_vector(to_unsigned( 83 , 8)),
                    5 => std_logic_vector(to_unsigned( 51 , 8)),
                    6 => std_logic_vector(to_unsigned( 3 , 8)),
                    7 => std_logic_vector(to_unsigned( 62 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1216 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 72, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 18 , 8)),
                    4 => std_logic_vector(to_unsigned( 83 , 8)),
                    5 => std_logic_vector(to_unsigned( 51 , 8)),
                    6 => std_logic_vector(to_unsigned( 3 , 8)),
                    7 => std_logic_vector(to_unsigned( 62 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1217 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 53, 8)),
                    1 => std_logic_vector(to_unsigned( 15 , 8)),
                    2 => std_logic_vector(to_unsigned( 116 , 8)),
                    3 => std_logic_vector(to_unsigned( 69 , 8)),
                    4 => std_logic_vector(to_unsigned( 83 , 8)),
                    5 => std_logic_vector(to_unsigned( 78 , 8)),
                    6 => std_logic_vector(to_unsigned( 7 , 8)),
                    7 => std_logic_vector(to_unsigned( 3 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1218 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),
                    1 => std_logic_vector(to_unsigned( 30 , 8)),
                    2 => std_logic_vector(to_unsigned( 60 , 8)),
                    3 => std_logic_vector(to_unsigned( 124 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 93 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1219 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),
                    1 => std_logic_vector(to_unsigned( 30 , 8)),
                    2 => std_logic_vector(to_unsigned( 60 , 8)),
                    3 => std_logic_vector(to_unsigned( 124 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 93 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1220 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 23 , 8)),
                    2 => std_logic_vector(to_unsigned( 27 , 8)),
                    3 => std_logic_vector(to_unsigned( 99 , 8)),
                    4 => std_logic_vector(to_unsigned( 51 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1221 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 66 , 8)),
                    2 => std_logic_vector(to_unsigned( 13 , 8)),
                    3 => std_logic_vector(to_unsigned( 73 , 8)),
                    4 => std_logic_vector(to_unsigned( 4 , 8)),
                    5 => std_logic_vector(to_unsigned( 38 , 8)),
                    6 => std_logic_vector(to_unsigned( 89 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1222 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 66 , 8)),
                    2 => std_logic_vector(to_unsigned( 13 , 8)),
                    3 => std_logic_vector(to_unsigned( 73 , 8)),
                    4 => std_logic_vector(to_unsigned( 4 , 8)),
                    5 => std_logic_vector(to_unsigned( 38 , 8)),
                    6 => std_logic_vector(to_unsigned( 89 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1223 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 45 , 8)),
                    3 => std_logic_vector(to_unsigned( 116 , 8)),
                    4 => std_logic_vector(to_unsigned( 12 , 8)),
                    5 => std_logic_vector(to_unsigned( 83 , 8)),
                    6 => std_logic_vector(to_unsigned( 56 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1224 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 94, 8)),
                    1 => std_logic_vector(to_unsigned( 65 , 8)),
                    2 => std_logic_vector(to_unsigned( 11 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 78 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 30 , 8)),
                    7 => std_logic_vector(to_unsigned( 116 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1225 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 94, 8)),
                    1 => std_logic_vector(to_unsigned( 65 , 8)),
                    2 => std_logic_vector(to_unsigned( 11 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 78 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 30 , 8)),
                    7 => std_logic_vector(to_unsigned( 116 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1226 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 33, 8)),
                    1 => std_logic_vector(to_unsigned( 20 , 8)),
                    2 => std_logic_vector(to_unsigned( 64 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 4 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 40 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1227 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 65, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 92 , 8)),
                    3 => std_logic_vector(to_unsigned( 12 , 8)),
                    4 => std_logic_vector(to_unsigned( 116 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 120 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1228 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 65, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 92 , 8)),
                    3 => std_logic_vector(to_unsigned( 12 , 8)),
                    4 => std_logic_vector(to_unsigned( 116 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 120 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1229 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 51, 8)),
                    1 => std_logic_vector(to_unsigned( 24 , 8)),
                    2 => std_logic_vector(to_unsigned( 93 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 117 , 8)),
                    6 => std_logic_vector(to_unsigned( 67 , 8)),
                    7 => std_logic_vector(to_unsigned( 105 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1230 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),
                    1 => std_logic_vector(to_unsigned( 38 , 8)),
                    2 => std_logic_vector(to_unsigned( 22 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 26 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 123 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1231 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),
                    1 => std_logic_vector(to_unsigned( 38 , 8)),
                    2 => std_logic_vector(to_unsigned( 22 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 26 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 123 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1232 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),
                    1 => std_logic_vector(to_unsigned( 38 , 8)),
                    2 => std_logic_vector(to_unsigned( 51 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 12 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 91 , 8)),
                    7 => std_logic_vector(to_unsigned( 121 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1233 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 54 , 8)),
                    2 => std_logic_vector(to_unsigned( 65 , 8)),
                    3 => std_logic_vector(to_unsigned( 109 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 29 , 8)),
                    6 => std_logic_vector(to_unsigned( 113 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1234 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 54 , 8)),
                    2 => std_logic_vector(to_unsigned( 65 , 8)),
                    3 => std_logic_vector(to_unsigned( 109 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 29 , 8)),
                    6 => std_logic_vector(to_unsigned( 113 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1235 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 45, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 36 , 8)),
                    4 => std_logic_vector(to_unsigned( 59 , 8)),
                    5 => std_logic_vector(to_unsigned( 18 , 8)),
                    6 => std_logic_vector(to_unsigned( 110 , 8)),
                    7 => std_logic_vector(to_unsigned( 0 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1236 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 37 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 120 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1237 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 87 , 8)),
                    2 => std_logic_vector(to_unsigned( 37 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 62 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 120 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1238 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 65, 8)),
                    1 => std_logic_vector(to_unsigned( 81 , 8)),
                    2 => std_logic_vector(to_unsigned( 18 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 76 , 8)),
                    5 => std_logic_vector(to_unsigned( 5 , 8)),
                    6 => std_logic_vector(to_unsigned( 60 , 8)),
                    7 => std_logic_vector(to_unsigned( 101 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1239 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),
                    1 => std_logic_vector(to_unsigned( 105 , 8)),
                    2 => std_logic_vector(to_unsigned( 75 , 8)),
                    3 => std_logic_vector(to_unsigned( 114 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 3 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1240 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),
                    1 => std_logic_vector(to_unsigned( 105 , 8)),
                    2 => std_logic_vector(to_unsigned( 75 , 8)),
                    3 => std_logic_vector(to_unsigned( 114 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 3 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1241 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 77 , 8)),
                    2 => std_logic_vector(to_unsigned( 6 , 8)),
                    3 => std_logic_vector(to_unsigned( 94 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 59 , 8)),
                    7 => std_logic_vector(to_unsigned( 105 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1242 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 90, 8)),
                    1 => std_logic_vector(to_unsigned( 115 , 8)),
                    2 => std_logic_vector(to_unsigned( 20 , 8)),
                    3 => std_logic_vector(to_unsigned( 11 , 8)),
                    4 => std_logic_vector(to_unsigned( 72 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 38 , 8)),
                    7 => std_logic_vector(to_unsigned( 53 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1243 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 90, 8)),
                    1 => std_logic_vector(to_unsigned( 115 , 8)),
                    2 => std_logic_vector(to_unsigned( 20 , 8)),
                    3 => std_logic_vector(to_unsigned( 11 , 8)),
                    4 => std_logic_vector(to_unsigned( 72 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 38 , 8)),
                    7 => std_logic_vector(to_unsigned( 53 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1244 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),
                    1 => std_logic_vector(to_unsigned( 68 , 8)),
                    2 => std_logic_vector(to_unsigned( 47 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 56 , 8)),
                    5 => std_logic_vector(to_unsigned( 94 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1245 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 54 , 8)),
                    2 => std_logic_vector(to_unsigned( 108 , 8)),
                    3 => std_logic_vector(to_unsigned( 39 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1246 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 54 , 8)),
                    2 => std_logic_vector(to_unsigned( 108 , 8)),
                    3 => std_logic_vector(to_unsigned( 39 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1247 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),
                    1 => std_logic_vector(to_unsigned( 42 , 8)),
                    2 => std_logic_vector(to_unsigned( 48 , 8)),
                    3 => std_logic_vector(to_unsigned( 123 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 116 , 8)),
                    6 => std_logic_vector(to_unsigned( 38 , 8)),
                    7 => std_logic_vector(to_unsigned( 108 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1248 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),
                    1 => std_logic_vector(to_unsigned( 57 , 8)),
                    2 => std_logic_vector(to_unsigned( 1 , 8)),
                    3 => std_logic_vector(to_unsigned( 17 , 8)),
                    4 => std_logic_vector(to_unsigned( 31 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 105 , 8)),
                    7 => std_logic_vector(to_unsigned( 38 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1249 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),
                    1 => std_logic_vector(to_unsigned( 57 , 8)),
                    2 => std_logic_vector(to_unsigned( 1 , 8)),
                    3 => std_logic_vector(to_unsigned( 17 , 8)),
                    4 => std_logic_vector(to_unsigned( 31 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 105 , 8)),
                    7 => std_logic_vector(to_unsigned( 38 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1250 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 106 , 8)),
                    2 => std_logic_vector(to_unsigned( 32 , 8)),
                    3 => std_logic_vector(to_unsigned( 0 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 92 , 8)),
                    6 => std_logic_vector(to_unsigned( 119 , 8)),
                    7 => std_logic_vector(to_unsigned( 9 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1251 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 112, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 63 , 8)),
                    3 => std_logic_vector(to_unsigned( 41 , 8)),
                    4 => std_logic_vector(to_unsigned( 21 , 8)),
                    5 => std_logic_vector(to_unsigned( 1 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 51 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1252 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 112, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 63 , 8)),
                    3 => std_logic_vector(to_unsigned( 41 , 8)),
                    4 => std_logic_vector(to_unsigned( 21 , 8)),
                    5 => std_logic_vector(to_unsigned( 1 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 51 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1253 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),
                    1 => std_logic_vector(to_unsigned( 82 , 8)),
                    2 => std_logic_vector(to_unsigned( 61 , 8)),
                    3 => std_logic_vector(to_unsigned( 5 , 8)),
                    4 => std_logic_vector(to_unsigned( 70 , 8)),
                    5 => std_logic_vector(to_unsigned( 18 , 8)),
                    6 => std_logic_vector(to_unsigned( 113 , 8)),
                    7 => std_logic_vector(to_unsigned( 105 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1254 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 20, 8)),
                    1 => std_logic_vector(to_unsigned( 7 , 8)),
                    2 => std_logic_vector(to_unsigned( 14 , 8)),
                    3 => std_logic_vector(to_unsigned( 25 , 8)),
                    4 => std_logic_vector(to_unsigned( 80 , 8)),
                    5 => std_logic_vector(to_unsigned( 52 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1255 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 20, 8)),
                    1 => std_logic_vector(to_unsigned( 7 , 8)),
                    2 => std_logic_vector(to_unsigned( 14 , 8)),
                    3 => std_logic_vector(to_unsigned( 25 , 8)),
                    4 => std_logic_vector(to_unsigned( 80 , 8)),
                    5 => std_logic_vector(to_unsigned( 52 , 8)),
                    6 => std_logic_vector(to_unsigned( 84 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1256 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 67, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 83 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 91 , 8)),
                    5 => std_logic_vector(to_unsigned( 15 , 8)),
                    6 => std_logic_vector(to_unsigned( 63 , 8)),
                    7 => std_logic_vector(to_unsigned( 118 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1257 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 90 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 64 , 8)),
                    5 => std_logic_vector(to_unsigned( 83 , 8)),
                    6 => std_logic_vector(to_unsigned( 117 , 8)),
                    7 => std_logic_vector(to_unsigned( 54 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1258 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 90 , 8)),
                    3 => std_logic_vector(to_unsigned( 32 , 8)),
                    4 => std_logic_vector(to_unsigned( 64 , 8)),
                    5 => std_logic_vector(to_unsigned( 83 , 8)),
                    6 => std_logic_vector(to_unsigned( 117 , 8)),
                    7 => std_logic_vector(to_unsigned( 54 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1259 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 30 , 8)),
                    2 => std_logic_vector(to_unsigned( 99 , 8)),
                    3 => std_logic_vector(to_unsigned( 123 , 8)),
                    4 => std_logic_vector(to_unsigned( 39 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 3 , 8)),
                    7 => std_logic_vector(to_unsigned( 56 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1260 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),
                    1 => std_logic_vector(to_unsigned( 67 , 8)),
                    2 => std_logic_vector(to_unsigned( 6 , 8)),
                    3 => std_logic_vector(to_unsigned( 10 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 45 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1261 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),
                    1 => std_logic_vector(to_unsigned( 67 , 8)),
                    2 => std_logic_vector(to_unsigned( 6 , 8)),
                    3 => std_logic_vector(to_unsigned( 10 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 45 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1262 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),
                    1 => std_logic_vector(to_unsigned( 58 , 8)),
                    2 => std_logic_vector(to_unsigned( 15 , 8)),
                    3 => std_logic_vector(to_unsigned( 54 , 8)),
                    4 => std_logic_vector(to_unsigned( 26 , 8)),
                    5 => std_logic_vector(to_unsigned( 73 , 8)),
                    6 => std_logic_vector(to_unsigned( 114 , 8)),
                    7 => std_logic_vector(to_unsigned( 20 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1263 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),
                    1 => std_logic_vector(to_unsigned( 84 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 50 , 8)),
                    4 => std_logic_vector(to_unsigned( 77 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 110 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1264 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),
                    1 => std_logic_vector(to_unsigned( 84 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 50 , 8)),
                    4 => std_logic_vector(to_unsigned( 77 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 110 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1265 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 37 , 8)),
                    2 => std_logic_vector(to_unsigned( 14 , 8)),
                    3 => std_logic_vector(to_unsigned( 98 , 8)),
                    4 => std_logic_vector(to_unsigned( 3 , 8)),
                    5 => std_logic_vector(to_unsigned( 30 , 8)),
                    6 => std_logic_vector(to_unsigned( 67 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1266 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 17 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 25 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 35 , 8)),
                    6 => std_logic_vector(to_unsigned( 123 , 8)),
                    7 => std_logic_vector(to_unsigned( 116 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1267 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 17 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 25 , 8)),
                    4 => std_logic_vector(to_unsigned( 58 , 8)),
                    5 => std_logic_vector(to_unsigned( 35 , 8)),
                    6 => std_logic_vector(to_unsigned( 123 , 8)),
                    7 => std_logic_vector(to_unsigned( 116 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1268 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 39, 8)),
                    1 => std_logic_vector(to_unsigned( 28 , 8)),
                    2 => std_logic_vector(to_unsigned( 54 , 8)),
                    3 => std_logic_vector(to_unsigned( 8 , 8)),
                    4 => std_logic_vector(to_unsigned( 43 , 8)),
                    5 => std_logic_vector(to_unsigned( 102 , 8)),
                    6 => std_logic_vector(to_unsigned( 82 , 8)),
                    7 => std_logic_vector(to_unsigned( 15 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1269 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),
                    1 => std_logic_vector(to_unsigned( 84 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 20 , 8)),
                    4 => std_logic_vector(to_unsigned( 70 , 8)),
                    5 => std_logic_vector(to_unsigned( 90 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 13 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1270 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),
                    1 => std_logic_vector(to_unsigned( 84 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 20 , 8)),
                    4 => std_logic_vector(to_unsigned( 70 , 8)),
                    5 => std_logic_vector(to_unsigned( 90 , 8)),
                    6 => std_logic_vector(to_unsigned( 62 , 8)),
                    7 => std_logic_vector(to_unsigned( 13 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1271 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 99, 8)),
                    1 => std_logic_vector(to_unsigned( 63 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 39 , 8)),
                    6 => std_logic_vector(to_unsigned( 56 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1272 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 2, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 117 , 8)),
                    3 => std_logic_vector(to_unsigned( 13 , 8)),
                    4 => std_logic_vector(to_unsigned( 21 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 38 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1273 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 2, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 117 , 8)),
                    3 => std_logic_vector(to_unsigned( 13 , 8)),
                    4 => std_logic_vector(to_unsigned( 21 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 38 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1274 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 92 , 8)),
                    3 => std_logic_vector(to_unsigned( 51 , 8)),
                    4 => std_logic_vector(to_unsigned( 84 , 8)),
                    5 => std_logic_vector(to_unsigned( 2 , 8)),
                    6 => std_logic_vector(to_unsigned( 14 , 8)),
                    7 => std_logic_vector(to_unsigned( 118 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1275 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 86 , 8)),
                    2 => std_logic_vector(to_unsigned( 104 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 37 , 8)),
                    6 => std_logic_vector(to_unsigned( 121 , 8)),
                    7 => std_logic_vector(to_unsigned( 67 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1276 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 86 , 8)),
                    2 => std_logic_vector(to_unsigned( 104 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 37 , 8)),
                    6 => std_logic_vector(to_unsigned( 121 , 8)),
                    7 => std_logic_vector(to_unsigned( 67 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1277 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 45, 8)),
                    1 => std_logic_vector(to_unsigned( 101 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 5 , 8)),
                    4 => std_logic_vector(to_unsigned( 90 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 68 , 8)),
                    7 => std_logic_vector(to_unsigned( 36 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1278 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 88 , 8)),
                    3 => std_logic_vector(to_unsigned( 11 , 8)),
                    4 => std_logic_vector(to_unsigned( 119 , 8)),
                    5 => std_logic_vector(to_unsigned( 56 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 97 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1279 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),
                    1 => std_logic_vector(to_unsigned( 78 , 8)),
                    2 => std_logic_vector(to_unsigned( 88 , 8)),
                    3 => std_logic_vector(to_unsigned( 11 , 8)),
                    4 => std_logic_vector(to_unsigned( 119 , 8)),
                    5 => std_logic_vector(to_unsigned( 56 , 8)),
                    6 => std_logic_vector(to_unsigned( 34 , 8)),
                    7 => std_logic_vector(to_unsigned( 97 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1280 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),
                    1 => std_logic_vector(to_unsigned( 43 , 8)),
                    2 => std_logic_vector(to_unsigned( 71 , 8)),
                    3 => std_logic_vector(to_unsigned( 49 , 8)),
                    4 => std_logic_vector(to_unsigned( 23 , 8)),
                    5 => std_logic_vector(to_unsigned( 27 , 8)),
                    6 => std_logic_vector(to_unsigned( 16 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1281 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 17, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 29 , 8)),
                    4 => std_logic_vector(to_unsigned( 50 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1282 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 17, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 107 , 8)),
                    3 => std_logic_vector(to_unsigned( 29 , 8)),
                    4 => std_logic_vector(to_unsigned( 50 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1283 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 72, 8)),
                    1 => std_logic_vector(to_unsigned( 91 , 8)),
                    2 => std_logic_vector(to_unsigned( 40 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 65 , 8)),
                    5 => std_logic_vector(to_unsigned( 77 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 26 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1284 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 48 , 8)),
                    3 => std_logic_vector(to_unsigned( 39 , 8)),
                    4 => std_logic_vector(to_unsigned( 11 , 8)),
                    5 => std_logic_vector(to_unsigned( 83 , 8)),
                    6 => std_logic_vector(to_unsigned( 117 , 8)),
                    7 => std_logic_vector(to_unsigned( 96 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1285 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 48 , 8)),
                    3 => std_logic_vector(to_unsigned( 39 , 8)),
                    4 => std_logic_vector(to_unsigned( 11 , 8)),
                    5 => std_logic_vector(to_unsigned( 83 , 8)),
                    6 => std_logic_vector(to_unsigned( 117 , 8)),
                    7 => std_logic_vector(to_unsigned( 96 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1286 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 77 , 8)),
                    2 => std_logic_vector(to_unsigned( 84 , 8)),
                    3 => std_logic_vector(to_unsigned( 53 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 109 , 8)),
                    6 => std_logic_vector(to_unsigned( 60 , 8)),
                    7 => std_logic_vector(to_unsigned( 23 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1287 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 6 , 8)),
                    2 => std_logic_vector(to_unsigned( 10 , 8)),
                    3 => std_logic_vector(to_unsigned( 111 , 8)),
                    4 => std_logic_vector(to_unsigned( 116 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 70 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1288 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 6 , 8)),
                    2 => std_logic_vector(to_unsigned( 10 , 8)),
                    3 => std_logic_vector(to_unsigned( 111 , 8)),
                    4 => std_logic_vector(to_unsigned( 116 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 70 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1289 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),
                    1 => std_logic_vector(to_unsigned( 81 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 85 , 8)),
                    4 => std_logic_vector(to_unsigned( 93 , 8)),
                    5 => std_logic_vector(to_unsigned( 68 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1290 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),
                    1 => std_logic_vector(to_unsigned( 51 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 36 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 68 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 60 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1291 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),
                    1 => std_logic_vector(to_unsigned( 51 , 8)),
                    2 => std_logic_vector(to_unsigned( 44 , 8)),
                    3 => std_logic_vector(to_unsigned( 36 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 68 , 8)),
                    6 => std_logic_vector(to_unsigned( 11 , 8)),
                    7 => std_logic_vector(to_unsigned( 60 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1292 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 58, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 114 , 8)),
                    3 => std_logic_vector(to_unsigned( 109 , 8)),
                    4 => std_logic_vector(to_unsigned( 24 , 8)),
                    5 => std_logic_vector(to_unsigned( 71 , 8)),
                    6 => std_logic_vector(to_unsigned( 77 , 8)),
                    7 => std_logic_vector(to_unsigned( 88 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1293 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 115 , 8)),
                    4 => std_logic_vector(to_unsigned( 122 , 8)),
                    5 => std_logic_vector(to_unsigned( 10 , 8)),
                    6 => std_logic_vector(to_unsigned( 50 , 8)),
                    7 => std_logic_vector(to_unsigned( 21 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1294 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 115 , 8)),
                    4 => std_logic_vector(to_unsigned( 122 , 8)),
                    5 => std_logic_vector(to_unsigned( 10 , 8)),
                    6 => std_logic_vector(to_unsigned( 50 , 8)),
                    7 => std_logic_vector(to_unsigned( 21 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1295 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 114, 8)),
                    1 => std_logic_vector(to_unsigned( 37 , 8)),
                    2 => std_logic_vector(to_unsigned( 18 , 8)),
                    3 => std_logic_vector(to_unsigned( 77 , 8)),
                    4 => std_logic_vector(to_unsigned( 52 , 8)),
                    5 => std_logic_vector(to_unsigned( 47 , 8)),
                    6 => std_logic_vector(to_unsigned( 120 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1296 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),
                    1 => std_logic_vector(to_unsigned( 46 , 8)),
                    2 => std_logic_vector(to_unsigned( 13 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 20 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1297 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),
                    1 => std_logic_vector(to_unsigned( 46 , 8)),
                    2 => std_logic_vector(to_unsigned( 13 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 20 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1298 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),
                    1 => std_logic_vector(to_unsigned( 59 , 8)),
                    2 => std_logic_vector(to_unsigned( 78 , 8)),
                    3 => std_logic_vector(to_unsigned( 5 , 8)),
                    4 => std_logic_vector(to_unsigned( 96 , 8)),
                    5 => std_logic_vector(to_unsigned( 118 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 33 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1299 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 96, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 19 , 8)),
                    3 => std_logic_vector(to_unsigned( 71 , 8)),
                    4 => std_logic_vector(to_unsigned( 92 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 110 , 8)),
                    7 => std_logic_vector(to_unsigned( 75 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1300 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 96, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 19 , 8)),
                    3 => std_logic_vector(to_unsigned( 71 , 8)),
                    4 => std_logic_vector(to_unsigned( 92 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 110 , 8)),
                    7 => std_logic_vector(to_unsigned( 75 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1301 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 62, 8)),
                    1 => std_logic_vector(to_unsigned( 72 , 8)),
                    2 => std_logic_vector(to_unsigned( 109 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 4 , 8)),
                    5 => std_logic_vector(to_unsigned( 17 , 8)),
                    6 => std_logic_vector(to_unsigned( 80 , 8)),
                    7 => std_logic_vector(to_unsigned( 94 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1302 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 40 , 8)),
                    3 => std_logic_vector(to_unsigned( 117 , 8)),
                    4 => std_logic_vector(to_unsigned( 103 , 8)),
                    5 => std_logic_vector(to_unsigned( 110 , 8)),
                    6 => std_logic_vector(to_unsigned( 56 , 8)),
                    7 => std_logic_vector(to_unsigned( 35 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1303 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 40 , 8)),
                    3 => std_logic_vector(to_unsigned( 117 , 8)),
                    4 => std_logic_vector(to_unsigned( 103 , 8)),
                    5 => std_logic_vector(to_unsigned( 110 , 8)),
                    6 => std_logic_vector(to_unsigned( 56 , 8)),
                    7 => std_logic_vector(to_unsigned( 35 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1304 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),
                    1 => std_logic_vector(to_unsigned( 95 , 8)),
                    2 => std_logic_vector(to_unsigned( 49 , 8)),
                    3 => std_logic_vector(to_unsigned( 115 , 8)),
                    4 => std_logic_vector(to_unsigned( 27 , 8)),
                    5 => std_logic_vector(to_unsigned( 108 , 8)),
                    6 => std_logic_vector(to_unsigned( 85 , 8)),
                    7 => std_logic_vector(to_unsigned( 70 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1305 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 23 , 8)),
                    2 => std_logic_vector(to_unsigned( 58 , 8)),
                    3 => std_logic_vector(to_unsigned( 96 , 8)),
                    4 => std_logic_vector(to_unsigned( 31 , 8)),
                    5 => std_logic_vector(to_unsigned( 120 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1306 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 23 , 8)),
                    2 => std_logic_vector(to_unsigned( 58 , 8)),
                    3 => std_logic_vector(to_unsigned( 96 , 8)),
                    4 => std_logic_vector(to_unsigned( 31 , 8)),
                    5 => std_logic_vector(to_unsigned( 120 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1307 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 58, 8)),
                    1 => std_logic_vector(to_unsigned( 66 , 8)),
                    2 => std_logic_vector(to_unsigned( 92 , 8)),
                    3 => std_logic_vector(to_unsigned( 78 , 8)),
                    4 => std_logic_vector(to_unsigned( 32 , 8)),
                    5 => std_logic_vector(to_unsigned( 7 , 8)),
                    6 => std_logic_vector(to_unsigned( 16 , 8)),
                    7 => std_logic_vector(to_unsigned( 104 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1308 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 9, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 115 , 8)),
                    3 => std_logic_vector(to_unsigned( 46 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 123 , 8)),
                    6 => std_logic_vector(to_unsigned( 78 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1309 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 9, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 115 , 8)),
                    3 => std_logic_vector(to_unsigned( 46 , 8)),
                    4 => std_logic_vector(to_unsigned( 100 , 8)),
                    5 => std_logic_vector(to_unsigned( 123 , 8)),
                    6 => std_logic_vector(to_unsigned( 78 , 8)),
                    7 => std_logic_vector(to_unsigned( 109 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1310 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 49 , 8)),
                    3 => std_logic_vector(to_unsigned( 106 , 8)),
                    4 => std_logic_vector(to_unsigned( 27 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 97 , 8)),
                    7 => std_logic_vector(to_unsigned( 40 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1311 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 9, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 59 , 8)),
                    4 => std_logic_vector(to_unsigned( 122 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 15 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1312 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 9, 8)),
                    1 => std_logic_vector(to_unsigned( 49 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 59 , 8)),
                    4 => std_logic_vector(to_unsigned( 122 , 8)),
                    5 => std_logic_vector(to_unsigned( 114 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 15 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1313 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),
                    1 => std_logic_vector(to_unsigned( 32 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 2 , 8)),
                    4 => std_logic_vector(to_unsigned( 121 , 8)),
                    5 => std_logic_vector(to_unsigned( 112 , 8)),
                    6 => std_logic_vector(to_unsigned( 26 , 8)),
                    7 => std_logic_vector(to_unsigned( 57 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1314 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 42 , 8)),
                    4 => std_logic_vector(to_unsigned( 1 , 8)),
                    5 => std_logic_vector(to_unsigned( 37 , 8)),
                    6 => std_logic_vector(to_unsigned( 77 , 8)),
                    7 => std_logic_vector(to_unsigned( 22 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1315 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 42 , 8)),
                    4 => std_logic_vector(to_unsigned( 1 , 8)),
                    5 => std_logic_vector(to_unsigned( 37 , 8)),
                    6 => std_logic_vector(to_unsigned( 77 , 8)),
                    7 => std_logic_vector(to_unsigned( 22 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1316 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),
                    1 => std_logic_vector(to_unsigned( 60 , 8)),
                    2 => std_logic_vector(to_unsigned( 80 , 8)),
                    3 => std_logic_vector(to_unsigned( 36 , 8)),
                    4 => std_logic_vector(to_unsigned( 96 , 8)),
                    5 => std_logic_vector(to_unsigned( 104 , 8)),
                    6 => std_logic_vector(to_unsigned( 6 , 8)),
                    7 => std_logic_vector(to_unsigned( 112 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1317 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 18 , 8)),
                    2 => std_logic_vector(to_unsigned( 68 , 8)),
                    3 => std_logic_vector(to_unsigned( 112 , 8)),
                    4 => std_logic_vector(to_unsigned( 9 , 8)),
                    5 => std_logic_vector(to_unsigned( 84 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 3 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1318 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 18 , 8)),
                    2 => std_logic_vector(to_unsigned( 68 , 8)),
                    3 => std_logic_vector(to_unsigned( 112 , 8)),
                    4 => std_logic_vector(to_unsigned( 9 , 8)),
                    5 => std_logic_vector(to_unsigned( 84 , 8)),
                    6 => std_logic_vector(to_unsigned( 99 , 8)),
                    7 => std_logic_vector(to_unsigned( 3 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1319 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),
                    1 => std_logic_vector(to_unsigned( 52 , 8)),
                    2 => std_logic_vector(to_unsigned( 28 , 8)),
                    3 => std_logic_vector(to_unsigned( 102 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 68 , 8)),
                    7 => std_logic_vector(to_unsigned( 47 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1320 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),
                    1 => std_logic_vector(to_unsigned( 29 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 49 , 8)),
                    6 => std_logic_vector(to_unsigned( 21 , 8)),
                    7 => std_logic_vector(to_unsigned( 54 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1321 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),
                    1 => std_logic_vector(to_unsigned( 29 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 49 , 8)),
                    6 => std_logic_vector(to_unsigned( 21 , 8)),
                    7 => std_logic_vector(to_unsigned( 54 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1322 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),
                    1 => std_logic_vector(to_unsigned( 112 , 8)),
                    2 => std_logic_vector(to_unsigned( 89 , 8)),
                    3 => std_logic_vector(to_unsigned( 67 , 8)),
                    4 => std_logic_vector(to_unsigned( 94 , 8)),
                    5 => std_logic_vector(to_unsigned( 118 , 8)),
                    6 => std_logic_vector(to_unsigned( 32 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1323 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 31 , 8)),
                    2 => std_logic_vector(to_unsigned( 50 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 67 , 8)),
                    5 => std_logic_vector(to_unsigned( 91 , 8)),
                    6 => std_logic_vector(to_unsigned( 25 , 8)),
                    7 => std_logic_vector(to_unsigned( 99 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1324 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),
                    1 => std_logic_vector(to_unsigned( 31 , 8)),
                    2 => std_logic_vector(to_unsigned( 50 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 67 , 8)),
                    5 => std_logic_vector(to_unsigned( 91 , 8)),
                    6 => std_logic_vector(to_unsigned( 25 , 8)),
                    7 => std_logic_vector(to_unsigned( 99 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1325 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),
                    1 => std_logic_vector(to_unsigned( 117 , 8)),
                    2 => std_logic_vector(to_unsigned( 51 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 10 , 8)),
                    6 => std_logic_vector(to_unsigned( 93 , 8)),
                    7 => std_logic_vector(to_unsigned( 41 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1326 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 9, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 104 , 8)),
                    3 => std_logic_vector(to_unsigned( 13 , 8)),
                    4 => std_logic_vector(to_unsigned( 55 , 8)),
                    5 => std_logic_vector(to_unsigned( 119 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1327 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 9, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 104 , 8)),
                    3 => std_logic_vector(to_unsigned( 13 , 8)),
                    4 => std_logic_vector(to_unsigned( 55 , 8)),
                    5 => std_logic_vector(to_unsigned( 119 , 8)),
                    6 => std_logic_vector(to_unsigned( 100 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1328 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 65, 8)),
                    1 => std_logic_vector(to_unsigned( 105 , 8)),
                    2 => std_logic_vector(to_unsigned( 42 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 88 , 8)),
                    6 => std_logic_vector(to_unsigned( 101 , 8)),
                    7 => std_logic_vector(to_unsigned( 69 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1329 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 45 , 8)),
                    2 => std_logic_vector(to_unsigned( 94 , 8)),
                    3 => std_logic_vector(to_unsigned( 37 , 8)),
                    4 => std_logic_vector(to_unsigned( 5 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 41 , 8)),
                    7 => std_logic_vector(to_unsigned( 67 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1330 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 45 , 8)),
                    2 => std_logic_vector(to_unsigned( 94 , 8)),
                    3 => std_logic_vector(to_unsigned( 37 , 8)),
                    4 => std_logic_vector(to_unsigned( 5 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 41 , 8)),
                    7 => std_logic_vector(to_unsigned( 67 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1331 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 67, 8)),
                    1 => std_logic_vector(to_unsigned( 53 , 8)),
                    2 => std_logic_vector(to_unsigned( 23 , 8)),
                    3 => std_logic_vector(to_unsigned( 60 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 15 , 8)),
                    6 => std_logic_vector(to_unsigned( 121 , 8)),
                    7 => std_logic_vector(to_unsigned( 108 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1332 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 88 , 8)),
                    3 => std_logic_vector(to_unsigned( 16 , 8)),
                    4 => std_logic_vector(to_unsigned( 2 , 8)),
                    5 => std_logic_vector(to_unsigned( 115 , 8)),
                    6 => std_logic_vector(to_unsigned( 26 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1333 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),
                    1 => std_logic_vector(to_unsigned( 122 , 8)),
                    2 => std_logic_vector(to_unsigned( 88 , 8)),
                    3 => std_logic_vector(to_unsigned( 16 , 8)),
                    4 => std_logic_vector(to_unsigned( 2 , 8)),
                    5 => std_logic_vector(to_unsigned( 115 , 8)),
                    6 => std_logic_vector(to_unsigned( 26 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1334 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 47, 8)),
                    1 => std_logic_vector(to_unsigned( 39 , 8)),
                    2 => std_logic_vector(to_unsigned( 102 , 8)),
                    3 => std_logic_vector(to_unsigned( 71 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 55 , 8)),
                    7 => std_logic_vector(to_unsigned( 75 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1335 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 85 , 8)),
                    2 => std_logic_vector(to_unsigned( 57 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 52 , 8)),
                    6 => std_logic_vector(to_unsigned( 10 , 8)),
                    7 => std_logic_vector(to_unsigned( 61 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1336 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),
                    1 => std_logic_vector(to_unsigned( 85 , 8)),
                    2 => std_logic_vector(to_unsigned( 57 , 8)),
                    3 => std_logic_vector(to_unsigned( 74 , 8)),
                    4 => std_logic_vector(to_unsigned( 95 , 8)),
                    5 => std_logic_vector(to_unsigned( 52 , 8)),
                    6 => std_logic_vector(to_unsigned( 10 , 8)),
                    7 => std_logic_vector(to_unsigned( 61 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1337 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),
                    1 => std_logic_vector(to_unsigned( 58 , 8)),
                    2 => std_logic_vector(to_unsigned( 42 , 8)),
                    3 => std_logic_vector(to_unsigned( 85 , 8)),
                    4 => std_logic_vector(to_unsigned( 37 , 8)),
                    5 => std_logic_vector(to_unsigned( 124 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1338 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 105, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 24 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 115 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1339 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 105, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 24 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 31 , 8)),
                    6 => std_logic_vector(to_unsigned( 115 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1340 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),
                    1 => std_logic_vector(to_unsigned( 111 , 8)),
                    2 => std_logic_vector(to_unsigned( 58 , 8)),
                    3 => std_logic_vector(to_unsigned( 11 , 8)),
                    4 => std_logic_vector(to_unsigned( 63 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 31 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1341 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 44 , 8)),
                    4 => std_logic_vector(to_unsigned( 19 , 8)),
                    5 => std_logic_vector(to_unsigned( 95 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1342 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),
                    1 => std_logic_vector(to_unsigned( 73 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 44 , 8)),
                    4 => std_logic_vector(to_unsigned( 19 , 8)),
                    5 => std_logic_vector(to_unsigned( 95 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1343 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),
                    1 => std_logic_vector(to_unsigned( 118 , 8)),
                    2 => std_logic_vector(to_unsigned( 50 , 8)),
                    3 => std_logic_vector(to_unsigned( 107 , 8)),
                    4 => std_logic_vector(to_unsigned( 77 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 60 , 8)),
                    7 => std_logic_vector(to_unsigned( 97 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1344 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),
                    1 => std_logic_vector(to_unsigned( 105 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 89 , 8)),
                    4 => std_logic_vector(to_unsigned( 53 , 8)),
                    5 => std_logic_vector(to_unsigned( 99 , 8)),
                    6 => std_logic_vector(to_unsigned( 45 , 8)),
                    7 => std_logic_vector(to_unsigned( 7 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1345 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),
                    1 => std_logic_vector(to_unsigned( 105 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 89 , 8)),
                    4 => std_logic_vector(to_unsigned( 53 , 8)),
                    5 => std_logic_vector(to_unsigned( 99 , 8)),
                    6 => std_logic_vector(to_unsigned( 45 , 8)),
                    7 => std_logic_vector(to_unsigned( 7 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1346 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),
                    1 => std_logic_vector(to_unsigned( 105 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 14 , 8)),
                    4 => std_logic_vector(to_unsigned( 70 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 42 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1347 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),
                    1 => std_logic_vector(to_unsigned( 52 , 8)),
                    2 => std_logic_vector(to_unsigned( 101 , 8)),
                    3 => std_logic_vector(to_unsigned( 77 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 33 , 8)),
                    6 => std_logic_vector(to_unsigned( 91 , 8)),
                    7 => std_logic_vector(to_unsigned( 40 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1348 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),
                    1 => std_logic_vector(to_unsigned( 52 , 8)),
                    2 => std_logic_vector(to_unsigned( 101 , 8)),
                    3 => std_logic_vector(to_unsigned( 77 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 33 , 8)),
                    6 => std_logic_vector(to_unsigned( 91 , 8)),
                    7 => std_logic_vector(to_unsigned( 40 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1349 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 114, 8)),
                    1 => std_logic_vector(to_unsigned( 5 , 8)),
                    2 => std_logic_vector(to_unsigned( 29 , 8)),
                    3 => std_logic_vector(to_unsigned( 40 , 8)),
                    4 => std_logic_vector(to_unsigned( 81 , 8)),
                    5 => std_logic_vector(to_unsigned( 118 , 8)),
                    6 => std_logic_vector(to_unsigned( 71 , 8)),
                    7 => std_logic_vector(to_unsigned( 91 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1350 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 38, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 108 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 60 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 54 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1351 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 38, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 108 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 60 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 54 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1352 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 118 , 8)),
                    3 => std_logic_vector(to_unsigned( 13 , 8)),
                    4 => std_logic_vector(to_unsigned( 24 , 8)),
                    5 => std_logic_vector(to_unsigned( 7 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 46 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1353 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),
                    1 => std_logic_vector(to_unsigned( 59 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 18 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 64 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 7 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1354 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),
                    1 => std_logic_vector(to_unsigned( 59 , 8)),
                    2 => std_logic_vector(to_unsigned( 55 , 8)),
                    3 => std_logic_vector(to_unsigned( 18 , 8)),
                    4 => std_logic_vector(to_unsigned( 35 , 8)),
                    5 => std_logic_vector(to_unsigned( 64 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 7 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1355 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 4, 8)),
                    1 => std_logic_vector(to_unsigned( 85 , 8)),
                    2 => std_logic_vector(to_unsigned( 103 , 8)),
                    3 => std_logic_vector(to_unsigned( 75 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 91 , 8)),
                    6 => std_logic_vector(to_unsigned( 25 , 8)),
                    7 => std_logic_vector(to_unsigned( 81 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1356 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 12, 8)),
                    1 => std_logic_vector(to_unsigned( 85 , 8)),
                    2 => std_logic_vector(to_unsigned( 96 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 2 , 8)),
                    5 => std_logic_vector(to_unsigned( 21 , 8)),
                    6 => std_logic_vector(to_unsigned( 79 , 8)),
                    7 => std_logic_vector(to_unsigned( 27 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1357 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 12, 8)),
                    1 => std_logic_vector(to_unsigned( 85 , 8)),
                    2 => std_logic_vector(to_unsigned( 96 , 8)),
                    3 => std_logic_vector(to_unsigned( 72 , 8)),
                    4 => std_logic_vector(to_unsigned( 2 , 8)),
                    5 => std_logic_vector(to_unsigned( 21 , 8)),
                    6 => std_logic_vector(to_unsigned( 79 , 8)),
                    7 => std_logic_vector(to_unsigned( 27 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1358 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 88 , 8)),
                    2 => std_logic_vector(to_unsigned( 67 , 8)),
                    3 => std_logic_vector(to_unsigned( 21 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 37 , 8)),
                    6 => std_logic_vector(to_unsigned( 44 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1359 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 32 , 8)),
                    3 => std_logic_vector(to_unsigned( 73 , 8)),
                    4 => std_logic_vector(to_unsigned( 4 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1360 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 32 , 8)),
                    3 => std_logic_vector(to_unsigned( 73 , 8)),
                    4 => std_logic_vector(to_unsigned( 4 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1361 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),
                    1 => std_logic_vector(to_unsigned( 109 , 8)),
                    2 => std_logic_vector(to_unsigned( 90 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 20 , 8)),
                    5 => std_logic_vector(to_unsigned( 28 , 8)),
                    6 => std_logic_vector(to_unsigned( 59 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1362 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 113 , 8)),
                    2 => std_logic_vector(to_unsigned( 43 , 8)),
                    3 => std_logic_vector(to_unsigned( 57 , 8)),
                    4 => std_logic_vector(to_unsigned( 123 , 8)),
                    5 => std_logic_vector(to_unsigned( 32 , 8)),
                    6 => std_logic_vector(to_unsigned( 85 , 8)),
                    7 => std_logic_vector(to_unsigned( 79 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1363 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),
                    1 => std_logic_vector(to_unsigned( 113 , 8)),
                    2 => std_logic_vector(to_unsigned( 43 , 8)),
                    3 => std_logic_vector(to_unsigned( 57 , 8)),
                    4 => std_logic_vector(to_unsigned( 123 , 8)),
                    5 => std_logic_vector(to_unsigned( 32 , 8)),
                    6 => std_logic_vector(to_unsigned( 85 , 8)),
                    7 => std_logic_vector(to_unsigned( 79 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1364 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 72, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 93 , 8)),
                    3 => std_logic_vector(to_unsigned( 103 , 8)),
                    4 => std_logic_vector(to_unsigned( 3 , 8)),
                    5 => std_logic_vector(to_unsigned( 39 , 8)),
                    6 => std_logic_vector(to_unsigned( 10 , 8)),
                    7 => std_logic_vector(to_unsigned( 45 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1365 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 18 , 8)),
                    3 => std_logic_vector(to_unsigned( 118 , 8)),
                    4 => std_logic_vector(to_unsigned( 80 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 43 , 8)),
                    7 => std_logic_vector(to_unsigned( 103 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1366 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 18 , 8)),
                    3 => std_logic_vector(to_unsigned( 118 , 8)),
                    4 => std_logic_vector(to_unsigned( 80 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 43 , 8)),
                    7 => std_logic_vector(to_unsigned( 103 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1367 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 16, 8)),
                    1 => std_logic_vector(to_unsigned( 32 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 69 , 8)),
                    5 => std_logic_vector(to_unsigned( 73 , 8)),
                    6 => std_logic_vector(to_unsigned( 107 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1368 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),
                    1 => std_logic_vector(to_unsigned( 33 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 18 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 4 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1369 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),
                    1 => std_logic_vector(to_unsigned( 33 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 18 , 8)),
                    4 => std_logic_vector(to_unsigned( 89 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 4 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1370 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 12 , 8)),
                    4 => std_logic_vector(to_unsigned( 107 , 8)),
                    5 => std_logic_vector(to_unsigned( 36 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 16 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1371 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 82 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 89 , 8)),
                    4 => std_logic_vector(to_unsigned( 98 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 109 , 8)),
                    7 => std_logic_vector(to_unsigned( 59 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1372 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),
                    1 => std_logic_vector(to_unsigned( 82 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 89 , 8)),
                    4 => std_logic_vector(to_unsigned( 98 , 8)),
                    5 => std_logic_vector(to_unsigned( 113 , 8)),
                    6 => std_logic_vector(to_unsigned( 109 , 8)),
                    7 => std_logic_vector(to_unsigned( 59 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1373 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 47, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 41 , 8)),
                    4 => std_logic_vector(to_unsigned( 2 , 8)),
                    5 => std_logic_vector(to_unsigned( 120 , 8)),
                    6 => std_logic_vector(to_unsigned( 79 , 8)),
                    7 => std_logic_vector(to_unsigned( 88 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1374 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 90, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 112 , 8)),
                    4 => std_logic_vector(to_unsigned( 6 , 8)),
                    5 => std_logic_vector(to_unsigned( 74 , 8)),
                    6 => std_logic_vector(to_unsigned( 16 , 8)),
                    7 => std_logic_vector(to_unsigned( 59 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1375 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 90, 8)),
                    1 => std_logic_vector(to_unsigned( 83 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 112 , 8)),
                    4 => std_logic_vector(to_unsigned( 6 , 8)),
                    5 => std_logic_vector(to_unsigned( 74 , 8)),
                    6 => std_logic_vector(to_unsigned( 16 , 8)),
                    7 => std_logic_vector(to_unsigned( 59 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1376 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 92 , 8)),
                    3 => std_logic_vector(to_unsigned( 50 , 8)),
                    4 => std_logic_vector(to_unsigned( 46 , 8)),
                    5 => std_logic_vector(to_unsigned( 117 , 8)),
                    6 => std_logic_vector(to_unsigned( 80 , 8)),
                    7 => std_logic_vector(to_unsigned( 56 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1377 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 96, 8)),
                    1 => std_logic_vector(to_unsigned( 60 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 42 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 26 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1378 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 96, 8)),
                    1 => std_logic_vector(to_unsigned( 60 , 8)),
                    2 => std_logic_vector(to_unsigned( 123 , 8)),
                    3 => std_logic_vector(to_unsigned( 42 , 8)),
                    4 => std_logic_vector(to_unsigned( 36 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 53 , 8)),
                    7 => std_logic_vector(to_unsigned( 26 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1379 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 5 , 8)),
                    2 => std_logic_vector(to_unsigned( 42 , 8)),
                    3 => std_logic_vector(to_unsigned( 33 , 8)),
                    4 => std_logic_vector(to_unsigned( 103 , 8)),
                    5 => std_logic_vector(to_unsigned( 116 , 8)),
                    6 => std_logic_vector(to_unsigned( 87 , 8)),
                    7 => std_logic_vector(to_unsigned( 58 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1380 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),
                    1 => std_logic_vector(to_unsigned( 63 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 106 , 8)),
                    5 => std_logic_vector(to_unsigned( 116 , 8)),
                    6 => std_logic_vector(to_unsigned( 77 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1381 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),
                    1 => std_logic_vector(to_unsigned( 63 , 8)),
                    2 => std_logic_vector(to_unsigned( 41 , 8)),
                    3 => std_logic_vector(to_unsigned( 47 , 8)),
                    4 => std_logic_vector(to_unsigned( 106 , 8)),
                    5 => std_logic_vector(to_unsigned( 116 , 8)),
                    6 => std_logic_vector(to_unsigned( 77 , 8)),
                    7 => std_logic_vector(to_unsigned( 95 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1382 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),
                    1 => std_logic_vector(to_unsigned( 5 , 8)),
                    2 => std_logic_vector(to_unsigned( 24 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 58 , 8)),
                    6 => std_logic_vector(to_unsigned( 87 , 8)),
                    7 => std_logic_vector(to_unsigned( 68 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1383 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),
                    1 => std_logic_vector(to_unsigned( 2 , 8)),
                    2 => std_logic_vector(to_unsigned( 11 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 116 , 8)),
                    6 => std_logic_vector(to_unsigned( 110 , 8)),
                    7 => std_logic_vector(to_unsigned( 96 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1384 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),
                    1 => std_logic_vector(to_unsigned( 2 , 8)),
                    2 => std_logic_vector(to_unsigned( 11 , 8)),
                    3 => std_logic_vector(to_unsigned( 30 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 116 , 8)),
                    6 => std_logic_vector(to_unsigned( 110 , 8)),
                    7 => std_logic_vector(to_unsigned( 96 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1385 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 114, 8)),
                    1 => std_logic_vector(to_unsigned( 66 , 8)),
                    2 => std_logic_vector(to_unsigned( 119 , 8)),
                    3 => std_logic_vector(to_unsigned( 13 , 8)),
                    4 => std_logic_vector(to_unsigned( 88 , 8)),
                    5 => std_logic_vector(to_unsigned( 78 , 8)),
                    6 => std_logic_vector(to_unsigned( 42 , 8)),
                    7 => std_logic_vector(to_unsigned( 73 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1386 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 115 , 8)),
                    3 => std_logic_vector(to_unsigned( 27 , 8)),
                    4 => std_logic_vector(to_unsigned( 119 , 8)),
                    5 => std_logic_vector(to_unsigned( 1 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1387 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 9 , 8)),
                    2 => std_logic_vector(to_unsigned( 115 , 8)),
                    3 => std_logic_vector(to_unsigned( 27 , 8)),
                    4 => std_logic_vector(to_unsigned( 119 , 8)),
                    5 => std_logic_vector(to_unsigned( 1 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1388 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),
                    1 => std_logic_vector(to_unsigned( 121 , 8)),
                    2 => std_logic_vector(to_unsigned( 54 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 9 , 8)),
                    5 => std_logic_vector(to_unsigned( 17 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 39 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1389 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 24 , 8)),
                    3 => std_logic_vector(to_unsigned( 120 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 101 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 40 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1390 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 116 , 8)),
                    2 => std_logic_vector(to_unsigned( 24 , 8)),
                    3 => std_logic_vector(to_unsigned( 120 , 8)),
                    4 => std_logic_vector(to_unsigned( 111 , 8)),
                    5 => std_logic_vector(to_unsigned( 101 , 8)),
                    6 => std_logic_vector(to_unsigned( 86 , 8)),
                    7 => std_logic_vector(to_unsigned( 40 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1391 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),
                    1 => std_logic_vector(to_unsigned( 24 , 8)),
                    2 => std_logic_vector(to_unsigned( 98 , 8)),
                    3 => std_logic_vector(to_unsigned( 76 , 8)),
                    4 => std_logic_vector(to_unsigned( 5 , 8)),
                    5 => std_logic_vector(to_unsigned( 36 , 8)),
                    6 => std_logic_vector(to_unsigned( 59 , 8)),
                    7 => std_logic_vector(to_unsigned( 11 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1392 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 71, 8)),
                    1 => std_logic_vector(to_unsigned( 85 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 93 , 8)),
                    4 => std_logic_vector(to_unsigned( 43 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 113 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1393 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 71, 8)),
                    1 => std_logic_vector(to_unsigned( 85 , 8)),
                    2 => std_logic_vector(to_unsigned( 7 , 8)),
                    3 => std_logic_vector(to_unsigned( 93 , 8)),
                    4 => std_logic_vector(to_unsigned( 43 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 113 , 8)),
                    7 => std_logic_vector(to_unsigned( 50 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1394 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 73, 8)),
                    1 => std_logic_vector(to_unsigned( 119 , 8)),
                    2 => std_logic_vector(to_unsigned( 99 , 8)),
                    3 => std_logic_vector(to_unsigned( 49 , 8)),
                    4 => std_logic_vector(to_unsigned( 44 , 8)),
                    5 => std_logic_vector(to_unsigned( 88 , 8)),
                    6 => std_logic_vector(to_unsigned( 115 , 8)),
                    7 => std_logic_vector(to_unsigned( 9 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1395 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 8 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 108 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 38 , 8)),
                    7 => std_logic_vector(to_unsigned( 32 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1396 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),
                    1 => std_logic_vector(to_unsigned( 8 , 8)),
                    2 => std_logic_vector(to_unsigned( 16 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 108 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 38 , 8)),
                    7 => std_logic_vector(to_unsigned( 32 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1397 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 117 , 8)),
                    2 => std_logic_vector(to_unsigned( 61 , 8)),
                    3 => std_logic_vector(to_unsigned( 88 , 8)),
                    4 => std_logic_vector(to_unsigned( 33 , 8)),
                    5 => std_logic_vector(to_unsigned( 100 , 8)),
                    6 => std_logic_vector(to_unsigned( 13 , 8)),
                    7 => std_logic_vector(to_unsigned( 112 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1398 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 58, 8)),
                    1 => std_logic_vector(to_unsigned( 100 , 8)),
                    2 => std_logic_vector(to_unsigned( 31 , 8)),
                    3 => std_logic_vector(to_unsigned( 109 , 8)),
                    4 => std_logic_vector(to_unsigned( 104 , 8)),
                    5 => std_logic_vector(to_unsigned( 20 , 8)),
                    6 => std_logic_vector(to_unsigned( 74 , 8)),
                    7 => std_logic_vector(to_unsigned( 11 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1399 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 58, 8)),
                    1 => std_logic_vector(to_unsigned( 100 , 8)),
                    2 => std_logic_vector(to_unsigned( 31 , 8)),
                    3 => std_logic_vector(to_unsigned( 109 , 8)),
                    4 => std_logic_vector(to_unsigned( 104 , 8)),
                    5 => std_logic_vector(to_unsigned( 20 , 8)),
                    6 => std_logic_vector(to_unsigned( 74 , 8)),
                    7 => std_logic_vector(to_unsigned( 11 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1400 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),
                    1 => std_logic_vector(to_unsigned( 70 , 8)),
                    2 => std_logic_vector(to_unsigned( 33 , 8)),
                    3 => std_logic_vector(to_unsigned( 77 , 8)),
                    4 => std_logic_vector(to_unsigned( 50 , 8)),
                    5 => std_logic_vector(to_unsigned( 61 , 8)),
                    6 => std_logic_vector(to_unsigned( 94 , 8)),
                    7 => std_logic_vector(to_unsigned( 46 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1401 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 37 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 44 , 8)),
                    4 => std_logic_vector(to_unsigned( 10 , 8)),
                    5 => std_logic_vector(to_unsigned( 2 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 108 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1402 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 37 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 44 , 8)),
                    4 => std_logic_vector(to_unsigned( 10 , 8)),
                    5 => std_logic_vector(to_unsigned( 2 , 8)),
                    6 => std_logic_vector(to_unsigned( 96 , 8)),
                    7 => std_logic_vector(to_unsigned( 108 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1403 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),
                    1 => std_logic_vector(to_unsigned( 92 , 8)),
                    2 => std_logic_vector(to_unsigned( 31 , 8)),
                    3 => std_logic_vector(to_unsigned( 118 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 84 , 8)),
                    6 => std_logic_vector(to_unsigned( 56 , 8)),
                    7 => std_logic_vector(to_unsigned( 1 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1404 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 71, 8)),
                    1 => std_logic_vector(to_unsigned( 119 , 8)),
                    2 => std_logic_vector(to_unsigned( 80 , 8)),
                    3 => std_logic_vector(to_unsigned( 49 , 8)),
                    4 => std_logic_vector(to_unsigned( 67 , 8)),
                    5 => std_logic_vector(to_unsigned( 32 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 14 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1405 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 71, 8)),
                    1 => std_logic_vector(to_unsigned( 119 , 8)),
                    2 => std_logic_vector(to_unsigned( 80 , 8)),
                    3 => std_logic_vector(to_unsigned( 49 , 8)),
                    4 => std_logic_vector(to_unsigned( 67 , 8)),
                    5 => std_logic_vector(to_unsigned( 32 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 14 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1406 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 4 , 8)),
                    2 => std_logic_vector(to_unsigned( 109 , 8)),
                    3 => std_logic_vector(to_unsigned( 14 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 82 , 8)),
                    6 => std_logic_vector(to_unsigned( 10 , 8)),
                    7 => std_logic_vector(to_unsigned( 71 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1407 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 81, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 27 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 2 , 8)),
                    6 => std_logic_vector(to_unsigned( 89 , 8)),
                    7 => std_logic_vector(to_unsigned( 121 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1408 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 81, 8)),
                    1 => std_logic_vector(to_unsigned( 69 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 27 , 8)),
                    4 => std_logic_vector(to_unsigned( 15 , 8)),
                    5 => std_logic_vector(to_unsigned( 2 , 8)),
                    6 => std_logic_vector(to_unsigned( 89 , 8)),
                    7 => std_logic_vector(to_unsigned( 121 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1409 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),
                    1 => std_logic_vector(to_unsigned( 96 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 70 , 8)),
                    4 => std_logic_vector(to_unsigned( 21 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 10 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1410 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 92 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 27 , 8)),
                    6 => std_logic_vector(to_unsigned( 88 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1411 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 124 , 8)),
                    3 => std_logic_vector(to_unsigned( 92 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 27 , 8)),
                    6 => std_logic_vector(to_unsigned( 88 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1412 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 93 , 8)),
                    3 => std_logic_vector(to_unsigned( 50 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 41 , 8)),
                    6 => std_logic_vector(to_unsigned( 63 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1413 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 20 , 8)),
                    2 => std_logic_vector(to_unsigned( 122 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 32 , 8)),
                    6 => std_logic_vector(to_unsigned( 67 , 8)),
                    7 => std_logic_vector(to_unsigned( 100 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1414 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 20 , 8)),
                    2 => std_logic_vector(to_unsigned( 122 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 71 , 8)),
                    5 => std_logic_vector(to_unsigned( 32 , 8)),
                    6 => std_logic_vector(to_unsigned( 67 , 8)),
                    7 => std_logic_vector(to_unsigned( 100 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1415 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 48 , 8)),
                    2 => std_logic_vector(to_unsigned( 102 , 8)),
                    3 => std_logic_vector(to_unsigned( 68 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 28 , 8)),
                    6 => std_logic_vector(to_unsigned( 95 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1416 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),
                    1 => std_logic_vector(to_unsigned( 12 , 8)),
                    2 => std_logic_vector(to_unsigned( 53 , 8)),
                    3 => std_logic_vector(to_unsigned( 60 , 8)),
                    4 => std_logic_vector(to_unsigned( 84 , 8)),
                    5 => std_logic_vector(to_unsigned( 38 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 16 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1417 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),
                    1 => std_logic_vector(to_unsigned( 12 , 8)),
                    2 => std_logic_vector(to_unsigned( 53 , 8)),
                    3 => std_logic_vector(to_unsigned( 60 , 8)),
                    4 => std_logic_vector(to_unsigned( 84 , 8)),
                    5 => std_logic_vector(to_unsigned( 38 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 16 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1418 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 92 , 8)),
                    3 => std_logic_vector(to_unsigned( 28 , 8)),
                    4 => std_logic_vector(to_unsigned( 65 , 8)),
                    5 => std_logic_vector(to_unsigned( 48 , 8)),
                    6 => std_logic_vector(to_unsigned( 111 , 8)),
                    7 => std_logic_vector(to_unsigned( 56 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1419 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),
                    1 => std_logic_vector(to_unsigned( 81 , 8)),
                    2 => std_logic_vector(to_unsigned( 115 , 8)),
                    3 => std_logic_vector(to_unsigned( 13 , 8)),
                    4 => std_logic_vector(to_unsigned( 25 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 104 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1420 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),
                    1 => std_logic_vector(to_unsigned( 81 , 8)),
                    2 => std_logic_vector(to_unsigned( 115 , 8)),
                    3 => std_logic_vector(to_unsigned( 13 , 8)),
                    4 => std_logic_vector(to_unsigned( 25 , 8)),
                    5 => std_logic_vector(to_unsigned( 9 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 104 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1421 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 3 , 8)),
                    3 => std_logic_vector(to_unsigned( 46 , 8)),
                    4 => std_logic_vector(to_unsigned( 16 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 66 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1422 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 18 , 8)),
                    4 => std_logic_vector(to_unsigned( 114 , 8)),
                    5 => std_logic_vector(to_unsigned( 23 , 8)),
                    6 => std_logic_vector(to_unsigned( 122 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1423 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),
                    1 => std_logic_vector(to_unsigned( 97 , 8)),
                    2 => std_logic_vector(to_unsigned( 8 , 8)),
                    3 => std_logic_vector(to_unsigned( 18 , 8)),
                    4 => std_logic_vector(to_unsigned( 114 , 8)),
                    5 => std_logic_vector(to_unsigned( 23 , 8)),
                    6 => std_logic_vector(to_unsigned( 122 , 8)),
                    7 => std_logic_vector(to_unsigned( 34 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1424 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 46, 8)),
                    1 => std_logic_vector(to_unsigned( 63 , 8)),
                    2 => std_logic_vector(to_unsigned( 99 , 8)),
                    3 => std_logic_vector(to_unsigned( 68 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 120 , 8)),
                    6 => std_logic_vector(to_unsigned( 59 , 8)),
                    7 => std_logic_vector(to_unsigned( 19 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1425 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 109 , 8)),
                    2 => std_logic_vector(to_unsigned( 91 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 68 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 113 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1426 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 109 , 8)),
                    2 => std_logic_vector(to_unsigned( 91 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 68 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 118 , 8)),
                    7 => std_logic_vector(to_unsigned( 113 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1427 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),
                    1 => std_logic_vector(to_unsigned( 34 , 8)),
                    2 => std_logic_vector(to_unsigned( 94 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 115 , 8)),
                    5 => std_logic_vector(to_unsigned( 66 , 8)),
                    6 => std_logic_vector(to_unsigned( 30 , 8)),
                    7 => std_logic_vector(to_unsigned( 83 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1428 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),
                    1 => std_logic_vector(to_unsigned( 46 , 8)),
                    2 => std_logic_vector(to_unsigned( 34 , 8)),
                    3 => std_logic_vector(to_unsigned( 114 , 8)),
                    4 => std_logic_vector(to_unsigned( 52 , 8)),
                    5 => std_logic_vector(to_unsigned( 14 , 8)),
                    6 => std_logic_vector(to_unsigned( 18 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1429 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),
                    1 => std_logic_vector(to_unsigned( 46 , 8)),
                    2 => std_logic_vector(to_unsigned( 34 , 8)),
                    3 => std_logic_vector(to_unsigned( 114 , 8)),
                    4 => std_logic_vector(to_unsigned( 52 , 8)),
                    5 => std_logic_vector(to_unsigned( 14 , 8)),
                    6 => std_logic_vector(to_unsigned( 18 , 8)),
                    7 => std_logic_vector(to_unsigned( 84 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1430 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 41, 8)),
                    1 => std_logic_vector(to_unsigned( 22 , 8)),
                    2 => std_logic_vector(to_unsigned( 87 , 8)),
                    3 => std_logic_vector(to_unsigned( 75 , 8)),
                    4 => std_logic_vector(to_unsigned( 106 , 8)),
                    5 => std_logic_vector(to_unsigned( 67 , 8)),
                    6 => std_logic_vector(to_unsigned( 9 , 8)),
                    7 => std_logic_vector(to_unsigned( 119 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1431 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 25 , 8)),
                    4 => std_logic_vector(to_unsigned( 40 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 8 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1432 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 110 , 8)),
                    3 => std_logic_vector(to_unsigned( 25 , 8)),
                    4 => std_logic_vector(to_unsigned( 40 , 8)),
                    5 => std_logic_vector(to_unsigned( 98 , 8)),
                    6 => std_logic_vector(to_unsigned( 8 , 8)),
                    7 => std_logic_vector(to_unsigned( 2 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1433 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),
                    1 => std_logic_vector(to_unsigned( 124 , 8)),
                    2 => std_logic_vector(to_unsigned( 75 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 9 , 8)),
                    5 => std_logic_vector(to_unsigned( 42 , 8)),
                    6 => std_logic_vector(to_unsigned( 28 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1434 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 106, 8)),
                    1 => std_logic_vector(to_unsigned( 64 , 8)),
                    2 => std_logic_vector(to_unsigned( 120 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 94 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1435 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 106, 8)),
                    1 => std_logic_vector(to_unsigned( 64 , 8)),
                    2 => std_logic_vector(to_unsigned( 120 , 8)),
                    3 => std_logic_vector(to_unsigned( 22 , 8)),
                    4 => std_logic_vector(to_unsigned( 29 , 8)),
                    5 => std_logic_vector(to_unsigned( 86 , 8)),
                    6 => std_logic_vector(to_unsigned( 47 , 8)),
                    7 => std_logic_vector(to_unsigned( 94 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1436 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 110, 8)),
                    1 => std_logic_vector(to_unsigned( 100 , 8)),
                    2 => std_logic_vector(to_unsigned( 37 , 8)),
                    3 => std_logic_vector(to_unsigned( 81 , 8)),
                    4 => std_logic_vector(to_unsigned( 30 , 8)),
                    5 => std_logic_vector(to_unsigned( 46 , 8)),
                    6 => std_logic_vector(to_unsigned( 74 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1437 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 51 , 8)),
                    2 => std_logic_vector(to_unsigned( 121 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 103 , 8)),
                    5 => std_logic_vector(to_unsigned( 92 , 8)),
                    6 => std_logic_vector(to_unsigned( 72 , 8)),
                    7 => std_logic_vector(to_unsigned( 8 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1438 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),
                    1 => std_logic_vector(to_unsigned( 51 , 8)),
                    2 => std_logic_vector(to_unsigned( 121 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 103 , 8)),
                    5 => std_logic_vector(to_unsigned( 92 , 8)),
                    6 => std_logic_vector(to_unsigned( 72 , 8)),
                    7 => std_logic_vector(to_unsigned( 8 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1439 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),
                    1 => std_logic_vector(to_unsigned( 60 , 8)),
                    2 => std_logic_vector(to_unsigned( 10 , 8)),
                    3 => std_logic_vector(to_unsigned( 15 , 8)),
                    4 => std_logic_vector(to_unsigned( 6 , 8)),
                    5 => std_logic_vector(to_unsigned( 79 , 8)),
                    6 => std_logic_vector(to_unsigned( 107 , 8)),
                    7 => std_logic_vector(to_unsigned( 21 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1440 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 45, 8)),
                    1 => std_logic_vector(to_unsigned( 52 , 8)),
                    2 => std_logic_vector(to_unsigned( 85 , 8)),
                    3 => std_logic_vector(to_unsigned( 12 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 117 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 67 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1441 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 45, 8)),
                    1 => std_logic_vector(to_unsigned( 52 , 8)),
                    2 => std_logic_vector(to_unsigned( 85 , 8)),
                    3 => std_logic_vector(to_unsigned( 12 , 8)),
                    4 => std_logic_vector(to_unsigned( 0 , 8)),
                    5 => std_logic_vector(to_unsigned( 117 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 67 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1442 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),
                    1 => std_logic_vector(to_unsigned( 121 , 8)),
                    2 => std_logic_vector(to_unsigned( 1 , 8)),
                    3 => std_logic_vector(to_unsigned( 8 , 8)),
                    4 => std_logic_vector(to_unsigned( 74 , 8)),
                    5 => std_logic_vector(to_unsigned( 12 , 8)),
                    6 => std_logic_vector(to_unsigned( 40 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1443 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 38, 8)),
                    1 => std_logic_vector(to_unsigned( 89 , 8)),
                    2 => std_logic_vector(to_unsigned( 6 , 8)),
                    3 => std_logic_vector(to_unsigned( 83 , 8)),
                    4 => std_logic_vector(to_unsigned( 94 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 26 , 8)),
                    7 => std_logic_vector(to_unsigned( 110 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1444 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 38, 8)),
                    1 => std_logic_vector(to_unsigned( 89 , 8)),
                    2 => std_logic_vector(to_unsigned( 6 , 8)),
                    3 => std_logic_vector(to_unsigned( 83 , 8)),
                    4 => std_logic_vector(to_unsigned( 94 , 8)),
                    5 => std_logic_vector(to_unsigned( 44 , 8)),
                    6 => std_logic_vector(to_unsigned( 26 , 8)),
                    7 => std_logic_vector(to_unsigned( 110 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1445 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),
                    1 => std_logic_vector(to_unsigned( 82 , 8)),
                    2 => std_logic_vector(to_unsigned( 36 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 40 , 8)),
                    5 => std_logic_vector(to_unsigned( 57 , 8)),
                    6 => std_logic_vector(to_unsigned( 74 , 8)),
                    7 => std_logic_vector(to_unsigned( 7 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1446 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 45 , 8)),
                    3 => std_logic_vector(to_unsigned( 15 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 94 , 8)),
                    6 => std_logic_vector(to_unsigned( 72 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1447 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),
                    1 => std_logic_vector(to_unsigned( 1 , 8)),
                    2 => std_logic_vector(to_unsigned( 45 , 8)),
                    3 => std_logic_vector(to_unsigned( 15 , 8)),
                    4 => std_logic_vector(to_unsigned( 112 , 8)),
                    5 => std_logic_vector(to_unsigned( 94 , 8)),
                    6 => std_logic_vector(to_unsigned( 72 , 8)),
                    7 => std_logic_vector(to_unsigned( 106 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1448 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 121, 8)),
                    1 => std_logic_vector(to_unsigned( 42 , 8)),
                    2 => std_logic_vector(to_unsigned( 79 , 8)),
                    3 => std_logic_vector(to_unsigned( 38 , 8)),
                    4 => std_logic_vector(to_unsigned( 92 , 8)),
                    5 => std_logic_vector(to_unsigned( 85 , 8)),
                    6 => std_logic_vector(to_unsigned( 28 , 8)),
                    7 => std_logic_vector(to_unsigned( 117 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1449 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 118 , 8)),
                    2 => std_logic_vector(to_unsigned( 84 , 8)),
                    3 => std_logic_vector(to_unsigned( 55 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 32 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1450 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 118 , 8)),
                    2 => std_logic_vector(to_unsigned( 84 , 8)),
                    3 => std_logic_vector(to_unsigned( 55 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 32 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 6 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1451 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),
                    1 => std_logic_vector(to_unsigned( 48 , 8)),
                    2 => std_logic_vector(to_unsigned( 17 , 8)),
                    3 => std_logic_vector(to_unsigned( 24 , 8)),
                    4 => std_logic_vector(to_unsigned( 61 , 8)),
                    5 => std_logic_vector(to_unsigned( 69 , 8)),
                    6 => std_logic_vector(to_unsigned( 2 , 8)),
                    7 => std_logic_vector(to_unsigned( 52 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1452 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 54, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 84 , 8)),
                    4 => std_logic_vector(to_unsigned( 45 , 8)),
                    5 => std_logic_vector(to_unsigned( 62 , 8)),
                    6 => std_logic_vector(to_unsigned( 72 , 8)),
                    7 => std_logic_vector(to_unsigned( 79 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1453 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 54, 8)),
                    1 => std_logic_vector(to_unsigned( 13 , 8)),
                    2 => std_logic_vector(to_unsigned( 5 , 8)),
                    3 => std_logic_vector(to_unsigned( 84 , 8)),
                    4 => std_logic_vector(to_unsigned( 45 , 8)),
                    5 => std_logic_vector(to_unsigned( 62 , 8)),
                    6 => std_logic_vector(to_unsigned( 72 , 8)),
                    7 => std_logic_vector(to_unsigned( 79 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1454 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 12, 8)),
                    1 => std_logic_vector(to_unsigned( 117 , 8)),
                    2 => std_logic_vector(to_unsigned( 3 , 8)),
                    3 => std_logic_vector(to_unsigned( 36 , 8)),
                    4 => std_logic_vector(to_unsigned( 69 , 8)),
                    5 => std_logic_vector(to_unsigned( 20 , 8)),
                    6 => std_logic_vector(to_unsigned( 108 , 8)),
                    7 => std_logic_vector(to_unsigned( 62 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1455 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 42, 8)),
                    1 => std_logic_vector(to_unsigned( 7 , 8)),
                    2 => std_logic_vector(to_unsigned( 29 , 8)),
                    3 => std_logic_vector(to_unsigned( 71 , 8)),
                    4 => std_logic_vector(to_unsigned( 103 , 8)),
                    5 => std_logic_vector(to_unsigned( 18 , 8)),
                    6 => std_logic_vector(to_unsigned( 1 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1456 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 42, 8)),
                    1 => std_logic_vector(to_unsigned( 7 , 8)),
                    2 => std_logic_vector(to_unsigned( 29 , 8)),
                    3 => std_logic_vector(to_unsigned( 71 , 8)),
                    4 => std_logic_vector(to_unsigned( 103 , 8)),
                    5 => std_logic_vector(to_unsigned( 18 , 8)),
                    6 => std_logic_vector(to_unsigned( 1 , 8)),
                    7 => std_logic_vector(to_unsigned( 86 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1457 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 64 , 8)),
                    2 => std_logic_vector(to_unsigned( 75 , 8)),
                    3 => std_logic_vector(to_unsigned( 1 , 8)),
                    4 => std_logic_vector(to_unsigned( 118 , 8)),
                    5 => std_logic_vector(to_unsigned( 89 , 8)),
                    6 => std_logic_vector(to_unsigned( 98 , 8)),
                    7 => std_logic_vector(to_unsigned( 80 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1458 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 124 , 8)),
                    2 => std_logic_vector(to_unsigned( 83 , 8)),
                    3 => std_logic_vector(to_unsigned( 23 , 8)),
                    4 => std_logic_vector(to_unsigned( 43 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 10 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1459 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),
                    1 => std_logic_vector(to_unsigned( 124 , 8)),
                    2 => std_logic_vector(to_unsigned( 83 , 8)),
                    3 => std_logic_vector(to_unsigned( 23 , 8)),
                    4 => std_logic_vector(to_unsigned( 43 , 8)),
                    5 => std_logic_vector(to_unsigned( 107 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 10 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1460 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),
                    1 => std_logic_vector(to_unsigned( 26 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 9 , 8)),
                    4 => std_logic_vector(to_unsigned( 86 , 8)),
                    5 => std_logic_vector(to_unsigned( 80 , 8)),
                    6 => std_logic_vector(to_unsigned( 105 , 8)),
                    7 => std_logic_vector(to_unsigned( 123 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1461 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 96, 8)),
                    1 => std_logic_vector(to_unsigned( 19 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 56 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 34 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 15 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1462 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 96, 8)),
                    1 => std_logic_vector(to_unsigned( 19 , 8)),
                    2 => std_logic_vector(to_unsigned( 77 , 8)),
                    3 => std_logic_vector(to_unsigned( 56 , 8)),
                    4 => std_logic_vector(to_unsigned( 109 , 8)),
                    5 => std_logic_vector(to_unsigned( 34 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 15 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1463 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 67, 8)),
                    1 => std_logic_vector(to_unsigned( 23 , 8)),
                    2 => std_logic_vector(to_unsigned( 102 , 8)),
                    3 => std_logic_vector(to_unsigned( 106 , 8)),
                    4 => std_logic_vector(to_unsigned( 72 , 8)),
                    5 => std_logic_vector(to_unsigned( 81 , 8)),
                    6 => std_logic_vector(to_unsigned( 2 , 8)),
                    7 => std_logic_vector(to_unsigned( 37 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1464 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 17 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 61 , 8)),
                    7 => std_logic_vector(to_unsigned( 48 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1465 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),
                    1 => std_logic_vector(to_unsigned( 55 , 8)),
                    2 => std_logic_vector(to_unsigned( 76 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 17 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 61 , 8)),
                    7 => std_logic_vector(to_unsigned( 48 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1466 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),
                    1 => std_logic_vector(to_unsigned( 58 , 8)),
                    2 => std_logic_vector(to_unsigned( 72 , 8)),
                    3 => std_logic_vector(to_unsigned( 48 , 8)),
                    4 => std_logic_vector(to_unsigned( 42 , 8)),
                    5 => std_logic_vector(to_unsigned( 112 , 8)),
                    6 => std_logic_vector(to_unsigned( 26 , 8)),
                    7 => std_logic_vector(to_unsigned( 52 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1467 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 53, 8)),
                    1 => std_logic_vector(to_unsigned( 107 , 8)),
                    2 => std_logic_vector(to_unsigned( 81 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 91 , 8)),
                    5 => std_logic_vector(to_unsigned( 49 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 13 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1468 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 53, 8)),
                    1 => std_logic_vector(to_unsigned( 107 , 8)),
                    2 => std_logic_vector(to_unsigned( 81 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 91 , 8)),
                    5 => std_logic_vector(to_unsigned( 49 , 8)),
                    6 => std_logic_vector(to_unsigned( 103 , 8)),
                    7 => std_logic_vector(to_unsigned( 13 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1469 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 4 , 8)),
                    3 => std_logic_vector(to_unsigned( 33 , 8)),
                    4 => std_logic_vector(to_unsigned( 49 , 8)),
                    5 => std_logic_vector(to_unsigned( 103 , 8)),
                    6 => std_logic_vector(to_unsigned( 0 , 8)),
                    7 => std_logic_vector(to_unsigned( 54 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1470 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 113 , 8)),
                    2 => std_logic_vector(to_unsigned( 9 , 8)),
                    3 => std_logic_vector(to_unsigned( 82 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 24 , 8)),
                    7 => std_logic_vector(to_unsigned( 88 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1471 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),
                    1 => std_logic_vector(to_unsigned( 113 , 8)),
                    2 => std_logic_vector(to_unsigned( 9 , 8)),
                    3 => std_logic_vector(to_unsigned( 82 , 8)),
                    4 => std_logic_vector(to_unsigned( 28 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 24 , 8)),
                    7 => std_logic_vector(to_unsigned( 88 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1472 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 15 , 8)),
                    2 => std_logic_vector(to_unsigned( 29 , 8)),
                    3 => std_logic_vector(to_unsigned( 79 , 8)),
                    4 => std_logic_vector(to_unsigned( 20 , 8)),
                    5 => std_logic_vector(to_unsigned( 106 , 8)),
                    6 => std_logic_vector(to_unsigned( 37 , 8)),
                    7 => std_logic_vector(to_unsigned( 85 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1473 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 72, 8)),
                    1 => std_logic_vector(to_unsigned( 50 , 8)),
                    2 => std_logic_vector(to_unsigned( 93 , 8)),
                    3 => std_logic_vector(to_unsigned( 84 , 8)),
                    4 => std_logic_vector(to_unsigned( 98 , 8)),
                    5 => std_logic_vector(to_unsigned( 88 , 8)),
                    6 => std_logic_vector(to_unsigned( 80 , 8)),
                    7 => std_logic_vector(to_unsigned( 35 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1474 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 72, 8)),
                    1 => std_logic_vector(to_unsigned( 50 , 8)),
                    2 => std_logic_vector(to_unsigned( 93 , 8)),
                    3 => std_logic_vector(to_unsigned( 84 , 8)),
                    4 => std_logic_vector(to_unsigned( 98 , 8)),
                    5 => std_logic_vector(to_unsigned( 88 , 8)),
                    6 => std_logic_vector(to_unsigned( 80 , 8)),
                    7 => std_logic_vector(to_unsigned( 35 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1475 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 118, 8)),
                    1 => std_logic_vector(to_unsigned( 36 , 8)),
                    2 => std_logic_vector(to_unsigned( 84 , 8)),
                    3 => std_logic_vector(to_unsigned( 52 , 8)),
                    4 => std_logic_vector(to_unsigned( 75 , 8)),
                    5 => std_logic_vector(to_unsigned( 70 , 8)),
                    6 => std_logic_vector(to_unsigned( 22 , 8)),
                    7 => std_logic_vector(to_unsigned( 102 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1476 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),
                    1 => std_logic_vector(to_unsigned( 62 , 8)),
                    2 => std_logic_vector(to_unsigned( 57 , 8)),
                    3 => std_logic_vector(to_unsigned( 83 , 8)),
                    4 => std_logic_vector(to_unsigned( 20 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 104 , 8)),
                    7 => std_logic_vector(to_unsigned( 51 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1477 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),
                    1 => std_logic_vector(to_unsigned( 62 , 8)),
                    2 => std_logic_vector(to_unsigned( 57 , 8)),
                    3 => std_logic_vector(to_unsigned( 83 , 8)),
                    4 => std_logic_vector(to_unsigned( 20 , 8)),
                    5 => std_logic_vector(to_unsigned( 26 , 8)),
                    6 => std_logic_vector(to_unsigned( 104 , 8)),
                    7 => std_logic_vector(to_unsigned( 51 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1478 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),
                    1 => std_logic_vector(to_unsigned( 25 , 8)),
                    2 => std_logic_vector(to_unsigned( 113 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 33 , 8)),
                    5 => std_logic_vector(to_unsigned( 119 , 8)),
                    6 => std_logic_vector(to_unsigned( 97 , 8)),
                    7 => std_logic_vector(to_unsigned( 47 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1479 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 113, 8)),
                    1 => std_logic_vector(to_unsigned( 7 , 8)),
                    2 => std_logic_vector(to_unsigned( 52 , 8)),
                    3 => std_logic_vector(to_unsigned( 122 , 8)),
                    4 => std_logic_vector(to_unsigned( 82 , 8)),
                    5 => std_logic_vector(to_unsigned( 64 , 8)),
                    6 => std_logic_vector(to_unsigned( 23 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1480 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 113, 8)),
                    1 => std_logic_vector(to_unsigned( 7 , 8)),
                    2 => std_logic_vector(to_unsigned( 52 , 8)),
                    3 => std_logic_vector(to_unsigned( 122 , 8)),
                    4 => std_logic_vector(to_unsigned( 82 , 8)),
                    5 => std_logic_vector(to_unsigned( 64 , 8)),
                    6 => std_logic_vector(to_unsigned( 23 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1481 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),
                    1 => std_logic_vector(to_unsigned( 32 , 8)),
                    2 => std_logic_vector(to_unsigned( 39 , 8)),
                    3 => std_logic_vector(to_unsigned( 80 , 8)),
                    4 => std_logic_vector(to_unsigned( 19 , 8)),
                    5 => std_logic_vector(to_unsigned( 97 , 8)),
                    6 => std_logic_vector(to_unsigned( 4 , 8)),
                    7 => std_logic_vector(to_unsigned( 74 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1482 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 25, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 59 , 8)),
                    3 => std_logic_vector(to_unsigned( 123 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 45 , 8)),
                    6 => std_logic_vector(to_unsigned( 64 , 8)),
                    7 => std_logic_vector(to_unsigned( 110 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1483 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 25, 8)),
                    1 => std_logic_vector(to_unsigned( 41 , 8)),
                    2 => std_logic_vector(to_unsigned( 59 , 8)),
                    3 => std_logic_vector(to_unsigned( 123 , 8)),
                    4 => std_logic_vector(to_unsigned( 102 , 8)),
                    5 => std_logic_vector(to_unsigned( 45 , 8)),
                    6 => std_logic_vector(to_unsigned( 64 , 8)),
                    7 => std_logic_vector(to_unsigned( 110 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1484 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),
                    1 => std_logic_vector(to_unsigned( 19 , 8)),
                    2 => std_logic_vector(to_unsigned( 54 , 8)),
                    3 => std_logic_vector(to_unsigned( 4 , 8)),
                    4 => std_logic_vector(to_unsigned( 113 , 8)),
                    5 => std_logic_vector(to_unsigned( 121 , 8)),
                    6 => std_logic_vector(to_unsigned( 80 , 8)),
                    7 => std_logic_vector(to_unsigned( 93 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1485 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 34 , 8)),
                    2 => std_logic_vector(to_unsigned( 58 , 8)),
                    3 => std_logic_vector(to_unsigned( 63 , 8)),
                    4 => std_logic_vector(to_unsigned( 11 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 2 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1486 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 34 , 8)),
                    2 => std_logic_vector(to_unsigned( 58 , 8)),
                    3 => std_logic_vector(to_unsigned( 63 , 8)),
                    4 => std_logic_vector(to_unsigned( 11 , 8)),
                    5 => std_logic_vector(to_unsigned( 16 , 8)),
                    6 => std_logic_vector(to_unsigned( 2 , 8)),
                    7 => std_logic_vector(to_unsigned( 89 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1487 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 40, 8)),
                    1 => std_logic_vector(to_unsigned( 104 , 8)),
                    2 => std_logic_vector(to_unsigned( 89 , 8)),
                    3 => std_logic_vector(to_unsigned( 34 , 8)),
                    4 => std_logic_vector(to_unsigned( 7 , 8)),
                    5 => std_logic_vector(to_unsigned( 22 , 8)),
                    6 => std_logic_vector(to_unsigned( 17 , 8)),
                    7 => std_logic_vector(to_unsigned( 72 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1488 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 33, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 94 , 8)),
                    3 => std_logic_vector(to_unsigned( 118 , 8)),
                    4 => std_logic_vector(to_unsigned( 106 , 8)),
                    5 => std_logic_vector(to_unsigned( 77 , 8)),
                    6 => std_logic_vector(to_unsigned( 58 , 8)),
                    7 => std_logic_vector(to_unsigned( 27 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1489 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 33, 8)),
                    1 => std_logic_vector(to_unsigned( 11 , 8)),
                    2 => std_logic_vector(to_unsigned( 94 , 8)),
                    3 => std_logic_vector(to_unsigned( 118 , 8)),
                    4 => std_logic_vector(to_unsigned( 106 , 8)),
                    5 => std_logic_vector(to_unsigned( 77 , 8)),
                    6 => std_logic_vector(to_unsigned( 58 , 8)),
                    7 => std_logic_vector(to_unsigned( 27 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1490 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),
                    1 => std_logic_vector(to_unsigned( 46 , 8)),
                    2 => std_logic_vector(to_unsigned( 3 , 8)),
                    3 => std_logic_vector(to_unsigned( 76 , 8)),
                    4 => std_logic_vector(to_unsigned( 52 , 8)),
                    5 => std_logic_vector(to_unsigned( 61 , 8)),
                    6 => std_logic_vector(to_unsigned( 41 , 8)),
                    7 => std_logic_vector(to_unsigned( 103 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1491 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 56 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 62 , 8)),
                    4 => std_logic_vector(to_unsigned( 1 , 8)),
                    5 => std_logic_vector(to_unsigned( 119 , 8)),
                    6 => std_logic_vector(to_unsigned( 114 , 8)),
                    7 => std_logic_vector(to_unsigned( 7 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1492 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),
                    1 => std_logic_vector(to_unsigned( 56 , 8)),
                    2 => std_logic_vector(to_unsigned( 95 , 8)),
                    3 => std_logic_vector(to_unsigned( 62 , 8)),
                    4 => std_logic_vector(to_unsigned( 1 , 8)),
                    5 => std_logic_vector(to_unsigned( 119 , 8)),
                    6 => std_logic_vector(to_unsigned( 114 , 8)),
                    7 => std_logic_vector(to_unsigned( 7 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1493 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),
                    1 => std_logic_vector(to_unsigned( 74 , 8)),
                    2 => std_logic_vector(to_unsigned( 66 , 8)),
                    3 => std_logic_vector(to_unsigned( 104 , 8)),
                    4 => std_logic_vector(to_unsigned( 52 , 8)),
                    5 => std_logic_vector(to_unsigned( 111 , 8)),
                    6 => std_logic_vector(to_unsigned( 39 , 8)),
                    7 => std_logic_vector(to_unsigned( 22 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1494 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),
                    1 => std_logic_vector(to_unsigned( 25 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 50 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 21 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1495 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),
                    1 => std_logic_vector(to_unsigned( 25 , 8)),
                    2 => std_logic_vector(to_unsigned( 0 , 8)),
                    3 => std_logic_vector(to_unsigned( 90 , 8)),
                    4 => std_logic_vector(to_unsigned( 50 , 8)),
                    5 => std_logic_vector(to_unsigned( 40 , 8)),
                    6 => std_logic_vector(to_unsigned( 21 , 8)),
                    7 => std_logic_vector(to_unsigned( 124 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1496 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 65, 8)),
                    1 => std_logic_vector(to_unsigned( 102 , 8)),
                    2 => std_logic_vector(to_unsigned( 34 , 8)),
                    3 => std_logic_vector(to_unsigned( 53 , 8)),
                    4 => std_logic_vector(to_unsigned( 124 , 8)),
                    5 => std_logic_vector(to_unsigned( 13 , 8)),
                    6 => std_logic_vector(to_unsigned( 19 , 8)),
                    7 => std_logic_vector(to_unsigned( 70 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1497 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),
                    1 => std_logic_vector(to_unsigned( 32 , 8)),
                    2 => std_logic_vector(to_unsigned( 101 , 8)),
                    3 => std_logic_vector(to_unsigned( 55 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 93 , 8)),
                    6 => std_logic_vector(to_unsigned( 2 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1498 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),
                    1 => std_logic_vector(to_unsigned( 32 , 8)),
                    2 => std_logic_vector(to_unsigned( 101 , 8)),
                    3 => std_logic_vector(to_unsigned( 55 , 8)),
                    4 => std_logic_vector(to_unsigned( 117 , 8)),
                    5 => std_logic_vector(to_unsigned( 93 , 8)),
                    6 => std_logic_vector(to_unsigned( 2 , 8)),
                    7 => std_logic_vector(to_unsigned( 63 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
         if i=1499 and is_next=1 then
            RAM <= (0 => std_logic_vector(to_unsigned( 16, 8)),
                    1 => std_logic_vector(to_unsigned( 65 , 8)),
                    2 => std_logic_vector(to_unsigned( 26 , 8)),
                    3 => std_logic_vector(to_unsigned( 59 , 8)),
                    4 => std_logic_vector(to_unsigned( 96 , 8)),
                    5 => std_logic_vector(to_unsigned( 105 , 8)),
                    6 => std_logic_vector(to_unsigned( 75 , 8)),
                    7 => std_logic_vector(to_unsigned( 49 , 8)),
                    8 => std_logic_vector(to_unsigned( addrs(i) , 8)),
        others => (others =>'0'));
    end if;
    
    end if;
end process;



test : process is
begin
if i < 1500 then
    wait for 100 ns;
    wait for c_CLOCK_PERIOD;
    tb_rst <= '1';
    wait for c_CLOCK_PERIOD;
    tb_rst <= '0';
    wait for c_CLOCK_PERIOD;
    tb_start <= '1';
    wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';

    -- Maschera di output = 0 - 129
    assert RAM(9) = std_logic_vector(to_unsigned( enc_addrs(i) , 8)) report "TEST FALLITO. Expected " & integer'image(enc_addrs(i)) & " found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

    i := i+1;
    is_next := 1;

    wait for c_CLOCK_PERIOD;
    wait for c_CLOCK_PERIOD;

    is_next := 0;

    if i=1500 then
        assert false report "Simulation Ended!, TEST PASSATO" severity failure;
    end if;
end if;
end process test;

end projecttb;




